

module vgg11
(
  input CLK,
  input RESETN,
  output reg irq,
  output reg [32-1:0] maxi_awaddr,
  output reg [8-1:0] maxi_awlen,
  output [3-1:0] maxi_awsize,
  output [2-1:0] maxi_awburst,
  output [1-1:0] maxi_awlock,
  output [4-1:0] maxi_awcache,
  output [3-1:0] maxi_awprot,
  output [4-1:0] maxi_awqos,
  output [2-1:0] maxi_awuser,
  output reg maxi_awvalid,
  input maxi_awready,
  output [32-1:0] maxi_wdata,
  output [4-1:0] maxi_wstrb,
  output maxi_wlast,
  output maxi_wvalid,
  input maxi_wready,
  input [2-1:0] maxi_bresp,
  input maxi_bvalid,
  output maxi_bready,
  output reg [32-1:0] maxi_araddr,
  output reg [8-1:0] maxi_arlen,
  output [3-1:0] maxi_arsize,
  output [2-1:0] maxi_arburst,
  output [1-1:0] maxi_arlock,
  output [4-1:0] maxi_arcache,
  output [3-1:0] maxi_arprot,
  output [4-1:0] maxi_arqos,
  output [2-1:0] maxi_aruser,
  output reg maxi_arvalid,
  input maxi_arready,
  input [32-1:0] maxi_rdata,
  input [2-1:0] maxi_rresp,
  input maxi_rlast,
  input maxi_rvalid,
  output maxi_rready,
  input [32-1:0] saxi_awaddr,
  input [4-1:0] saxi_awcache,
  input [3-1:0] saxi_awprot,
  input saxi_awvalid,
  output saxi_awready,
  input [32-1:0] saxi_wdata,
  input [4-1:0] saxi_wstrb,
  input saxi_wvalid,
  output saxi_wready,
  output [2-1:0] saxi_bresp,
  output reg saxi_bvalid,
  input saxi_bready,
  input [32-1:0] saxi_araddr,
  input [4-1:0] saxi_arcache,
  input [3-1:0] saxi_arprot,
  input saxi_arvalid,
  output saxi_arready,
  output reg [32-1:0] saxi_rdata,
  output [2-1:0] saxi_rresp,
  output reg saxi_rvalid,
  input saxi_rready
);

  wire RESETN_inv;
  assign RESETN_inv = !RESETN;
  wire RESETN_inv_buf;
  reg _RESETN_inv_1;
  reg _RESETN_inv_2;
  assign RESETN_inv_buf = _RESETN_inv_2;
  assign maxi_awsize = 2;
  assign maxi_awburst = 1;
  assign maxi_awlock = 0;
  assign maxi_awcache = 3;
  assign maxi_awprot = 0;
  assign maxi_awqos = 0;
  assign maxi_awuser = 0;
  reg [32-1:0] _maxi_wdata_sb_0;
  reg [4-1:0] _maxi_wstrb_sb_0;
  reg _maxi_wlast_sb_0;
  reg _maxi_wvalid_sb_0;
  wire _maxi_wready_sb_0;
  wire _sb_maxi_writedata_s_value_0;
  assign _sb_maxi_writedata_s_value_0 = _maxi_wlast_sb_0;
  wire [4-1:0] _sb_maxi_writedata_s_value_1;
  assign _sb_maxi_writedata_s_value_1 = _maxi_wstrb_sb_0;
  wire [32-1:0] _sb_maxi_writedata_s_value_2;
  assign _sb_maxi_writedata_s_value_2 = _maxi_wdata_sb_0;
  wire [37-1:0] _sb_maxi_writedata_s_data_3;
  assign _sb_maxi_writedata_s_data_3 = { _sb_maxi_writedata_s_value_0, _sb_maxi_writedata_s_value_1, _sb_maxi_writedata_s_value_2 };
  wire _sb_maxi_writedata_s_valid_4;
  assign _sb_maxi_writedata_s_valid_4 = _maxi_wvalid_sb_0;
  wire _sb_maxi_writedata_m_ready_5;
  assign _sb_maxi_writedata_m_ready_5 = maxi_wready;
  reg [37-1:0] _sb_maxi_writedata_data_6;
  reg _sb_maxi_writedata_valid_7;
  wire _sb_maxi_writedata_ready_8;
  reg [37-1:0] _sb_maxi_writedata_tmp_data_9;
  reg _sb_maxi_writedata_tmp_valid_10;
  wire [37-1:0] _sb_maxi_writedata_next_data_11;
  wire _sb_maxi_writedata_next_valid_12;
  assign _sb_maxi_writedata_ready_8 = !_sb_maxi_writedata_tmp_valid_10;
  assign _sb_maxi_writedata_next_data_11 = (_sb_maxi_writedata_tmp_valid_10)? _sb_maxi_writedata_tmp_data_9 : _sb_maxi_writedata_s_data_3;
  assign _sb_maxi_writedata_next_valid_12 = _sb_maxi_writedata_tmp_valid_10 || _sb_maxi_writedata_s_valid_4;
  wire _sb_maxi_writedata_m_value_13;
  assign _sb_maxi_writedata_m_value_13 = _sb_maxi_writedata_data_6[36:36];
  wire [4-1:0] _sb_maxi_writedata_m_value_14;
  assign _sb_maxi_writedata_m_value_14 = _sb_maxi_writedata_data_6[35:32];
  wire [32-1:0] _sb_maxi_writedata_m_value_15;
  assign _sb_maxi_writedata_m_value_15 = _sb_maxi_writedata_data_6[31:0];
  assign _maxi_wready_sb_0 = _sb_maxi_writedata_ready_8;
  assign maxi_wdata = _sb_maxi_writedata_m_value_15;
  assign maxi_wstrb = _sb_maxi_writedata_m_value_14;
  assign maxi_wlast = _sb_maxi_writedata_m_value_13;
  assign maxi_wvalid = _sb_maxi_writedata_valid_7;
  assign maxi_bready = 1;
  assign maxi_arsize = 2;
  assign maxi_arburst = 1;
  assign maxi_arlock = 0;
  assign maxi_arcache = 3;
  assign maxi_arprot = 0;
  assign maxi_arqos = 0;
  assign maxi_aruser = 0;
  wire [32-1:0] _maxi_rdata_sb_0;
  wire _maxi_rlast_sb_0;
  wire _maxi_rvalid_sb_0;
  wire _maxi_rready_sb_0;
  wire _sb_maxi_readdata_s_value_16;
  assign _sb_maxi_readdata_s_value_16 = maxi_rlast;
  wire [32-1:0] _sb_maxi_readdata_s_value_17;
  assign _sb_maxi_readdata_s_value_17 = maxi_rdata;
  wire [33-1:0] _sb_maxi_readdata_s_data_18;
  assign _sb_maxi_readdata_s_data_18 = { _sb_maxi_readdata_s_value_16, _sb_maxi_readdata_s_value_17 };
  wire _sb_maxi_readdata_s_valid_19;
  assign _sb_maxi_readdata_s_valid_19 = maxi_rvalid;
  wire _sb_maxi_readdata_m_ready_20;
  assign _sb_maxi_readdata_m_ready_20 = _maxi_rready_sb_0;
  reg [33-1:0] _sb_maxi_readdata_data_21;
  reg _sb_maxi_readdata_valid_22;
  wire _sb_maxi_readdata_ready_23;
  reg [33-1:0] _sb_maxi_readdata_tmp_data_24;
  reg _sb_maxi_readdata_tmp_valid_25;
  wire [33-1:0] _sb_maxi_readdata_next_data_26;
  wire _sb_maxi_readdata_next_valid_27;
  assign _sb_maxi_readdata_ready_23 = !_sb_maxi_readdata_tmp_valid_25;
  assign _sb_maxi_readdata_next_data_26 = (_sb_maxi_readdata_tmp_valid_25)? _sb_maxi_readdata_tmp_data_24 : _sb_maxi_readdata_s_data_18;
  assign _sb_maxi_readdata_next_valid_27 = _sb_maxi_readdata_tmp_valid_25 || _sb_maxi_readdata_s_valid_19;
  wire _sb_maxi_readdata_m_value_28;
  assign _sb_maxi_readdata_m_value_28 = _sb_maxi_readdata_data_21[32:32];
  wire [32-1:0] _sb_maxi_readdata_m_value_29;
  assign _sb_maxi_readdata_m_value_29 = _sb_maxi_readdata_data_21[31:0];
  assign _maxi_rdata_sb_0 = _sb_maxi_readdata_m_value_29;
  assign _maxi_rlast_sb_0 = _sb_maxi_readdata_m_value_28;
  assign _maxi_rvalid_sb_0 = _sb_maxi_readdata_valid_22;
  assign maxi_rready = _sb_maxi_readdata_ready_23;
  reg [3-1:0] _maxi_outstanding_wcount;
  wire _maxi_has_outstanding_write;
  assign _maxi_has_outstanding_write = (_maxi_outstanding_wcount > 0) || maxi_awvalid;
  reg _maxi_read_start;
  reg [8-1:0] _maxi_read_op_sel;
  reg [32-1:0] _maxi_read_global_addr;
  reg [33-1:0] _maxi_read_global_size;
  reg [32-1:0] _maxi_read_local_addr;
  reg [32-1:0] _maxi_read_local_stride;
  reg [33-1:0] _maxi_read_local_size;
  reg [32-1:0] _maxi_read_local_blocksize;
  wire _maxi_read_req_fifo_enq;
  wire [137-1:0] _maxi_read_req_fifo_wdata;
  wire _maxi_read_req_fifo_full;
  wire _maxi_read_req_fifo_almost_full;
  wire _maxi_read_req_fifo_deq;
  wire [137-1:0] _maxi_read_req_fifo_rdata;
  wire _maxi_read_req_fifo_empty;
  wire _maxi_read_req_fifo_almost_empty;

  _maxi_read_req_fifo
  inst__maxi_read_req_fifo
  (
    .CLK(CLK),
    .RST(RESETN_inv_buf),
    ._maxi_read_req_fifo_enq(_maxi_read_req_fifo_enq),
    ._maxi_read_req_fifo_wdata(_maxi_read_req_fifo_wdata),
    ._maxi_read_req_fifo_full(_maxi_read_req_fifo_full),
    ._maxi_read_req_fifo_almost_full(_maxi_read_req_fifo_almost_full),
    ._maxi_read_req_fifo_deq(_maxi_read_req_fifo_deq),
    ._maxi_read_req_fifo_rdata(_maxi_read_req_fifo_rdata),
    ._maxi_read_req_fifo_empty(_maxi_read_req_fifo_empty),
    ._maxi_read_req_fifo_almost_empty(_maxi_read_req_fifo_almost_empty)
  );

  reg [4-1:0] count__maxi_read_req_fifo;
  wire [8-1:0] _maxi_read_op_sel_fifo;
  wire [32-1:0] _maxi_read_local_addr_fifo;
  wire [32-1:0] _maxi_read_local_stride_fifo;
  wire [33-1:0] _maxi_read_local_size_fifo;
  wire [32-1:0] _maxi_read_local_blocksize_fifo;
  wire [8-1:0] unpack_read_req_op_sel_30;
  wire [32-1:0] unpack_read_req_local_addr_31;
  wire [32-1:0] unpack_read_req_local_stride_32;
  wire [33-1:0] unpack_read_req_local_size_33;
  wire [32-1:0] unpack_read_req_local_blocksize_34;
  assign unpack_read_req_op_sel_30 = _maxi_read_req_fifo_rdata[136:129];
  assign unpack_read_req_local_addr_31 = _maxi_read_req_fifo_rdata[128:97];
  assign unpack_read_req_local_stride_32 = _maxi_read_req_fifo_rdata[96:65];
  assign unpack_read_req_local_size_33 = _maxi_read_req_fifo_rdata[64:32];
  assign unpack_read_req_local_blocksize_34 = _maxi_read_req_fifo_rdata[31:0];
  assign _maxi_read_op_sel_fifo = unpack_read_req_op_sel_30;
  assign _maxi_read_local_addr_fifo = unpack_read_req_local_addr_31;
  assign _maxi_read_local_stride_fifo = unpack_read_req_local_stride_32;
  assign _maxi_read_local_size_fifo = unpack_read_req_local_size_33;
  assign _maxi_read_local_blocksize_fifo = unpack_read_req_local_blocksize_34;
  reg [8-1:0] _maxi_read_op_sel_buf;
  reg [32-1:0] _maxi_read_local_addr_buf;
  reg [32-1:0] _maxi_read_local_stride_buf;
  reg [33-1:0] _maxi_read_local_size_buf;
  reg [32-1:0] _maxi_read_local_blocksize_buf;
  reg _maxi_read_req_busy;
  reg _maxi_read_data_busy;
  wire _maxi_read_req_idle;
  wire _maxi_read_data_idle;
  wire _maxi_read_idle;
  assign _maxi_read_req_idle = !_maxi_read_start && !_maxi_read_req_busy;
  assign _maxi_read_data_idle = _maxi_read_req_fifo_empty && !_maxi_read_data_busy;
  assign _maxi_read_idle = _maxi_read_req_idle && _maxi_read_data_idle;
  reg _maxi_write_start;
  reg [8-1:0] _maxi_write_op_sel;
  reg [32-1:0] _maxi_write_global_addr;
  reg [33-1:0] _maxi_write_global_size;
  reg [32-1:0] _maxi_write_local_addr;
  reg [32-1:0] _maxi_write_local_stride;
  reg [33-1:0] _maxi_write_local_size;
  reg [32-1:0] _maxi_write_local_blocksize;
  wire _maxi_write_req_fifo_enq;
  wire [137-1:0] _maxi_write_req_fifo_wdata;
  wire _maxi_write_req_fifo_full;
  wire _maxi_write_req_fifo_almost_full;
  wire _maxi_write_req_fifo_deq;
  wire [137-1:0] _maxi_write_req_fifo_rdata;
  wire _maxi_write_req_fifo_empty;
  wire _maxi_write_req_fifo_almost_empty;

  _maxi_write_req_fifo
  inst__maxi_write_req_fifo
  (
    .CLK(CLK),
    .RST(RESETN_inv_buf),
    ._maxi_write_req_fifo_enq(_maxi_write_req_fifo_enq),
    ._maxi_write_req_fifo_wdata(_maxi_write_req_fifo_wdata),
    ._maxi_write_req_fifo_full(_maxi_write_req_fifo_full),
    ._maxi_write_req_fifo_almost_full(_maxi_write_req_fifo_almost_full),
    ._maxi_write_req_fifo_deq(_maxi_write_req_fifo_deq),
    ._maxi_write_req_fifo_rdata(_maxi_write_req_fifo_rdata),
    ._maxi_write_req_fifo_empty(_maxi_write_req_fifo_empty),
    ._maxi_write_req_fifo_almost_empty(_maxi_write_req_fifo_almost_empty)
  );

  reg [4-1:0] count__maxi_write_req_fifo;
  wire [8-1:0] _maxi_write_op_sel_fifo;
  wire [32-1:0] _maxi_write_local_addr_fifo;
  wire [32-1:0] _maxi_write_local_stride_fifo;
  wire [33-1:0] _maxi_write_size_fifo;
  wire [32-1:0] _maxi_write_local_blocksize_fifo;
  wire [8-1:0] unpack_write_req_op_sel_35;
  wire [32-1:0] unpack_write_req_local_addr_36;
  wire [32-1:0] unpack_write_req_local_stride_37;
  wire [33-1:0] unpack_write_req_size_38;
  wire [32-1:0] unpack_write_req_local_blocksize_39;
  assign unpack_write_req_op_sel_35 = _maxi_write_req_fifo_rdata[136:129];
  assign unpack_write_req_local_addr_36 = _maxi_write_req_fifo_rdata[128:97];
  assign unpack_write_req_local_stride_37 = _maxi_write_req_fifo_rdata[96:65];
  assign unpack_write_req_size_38 = _maxi_write_req_fifo_rdata[64:32];
  assign unpack_write_req_local_blocksize_39 = _maxi_write_req_fifo_rdata[31:0];
  assign _maxi_write_op_sel_fifo = unpack_write_req_op_sel_35;
  assign _maxi_write_local_addr_fifo = unpack_write_req_local_addr_36;
  assign _maxi_write_local_stride_fifo = unpack_write_req_local_stride_37;
  assign _maxi_write_size_fifo = unpack_write_req_size_38;
  assign _maxi_write_local_blocksize_fifo = unpack_write_req_local_blocksize_39;
  reg [8-1:0] _maxi_write_op_sel_buf;
  reg [32-1:0] _maxi_write_local_addr_buf;
  reg [32-1:0] _maxi_write_local_stride_buf;
  reg [33-1:0] _maxi_write_size_buf;
  reg [32-1:0] _maxi_write_local_blocksize_buf;
  reg _maxi_write_req_busy;
  reg _maxi_write_data_busy;
  wire _maxi_write_req_idle;
  wire _maxi_write_data_idle;
  wire _maxi_write_idle;
  assign _maxi_write_req_idle = !_maxi_write_start && !_maxi_write_req_busy;
  assign _maxi_write_data_idle = _maxi_write_req_fifo_empty && !_maxi_write_data_busy;
  assign _maxi_write_idle = _maxi_write_req_idle && _maxi_write_data_idle;
  reg [32-1:0] _maxi_global_base_addr;
  assign saxi_bresp = 0;
  assign saxi_rresp = 0;
  reg signed [32-1:0] _saxi_register_0;
  reg signed [32-1:0] _saxi_register_1;
  reg signed [32-1:0] _saxi_register_2;
  reg signed [32-1:0] _saxi_register_3;
  reg signed [32-1:0] _saxi_register_4;
  reg signed [32-1:0] _saxi_register_5;
  reg signed [32-1:0] _saxi_register_6;
  reg signed [32-1:0] _saxi_register_7;
  reg signed [32-1:0] _saxi_register_8;
  reg signed [32-1:0] _saxi_register_9;
  reg signed [32-1:0] _saxi_register_10;
  reg signed [32-1:0] _saxi_register_11;
  reg signed [32-1:0] _saxi_register_12;
  reg signed [32-1:0] _saxi_register_13;
  reg signed [32-1:0] _saxi_register_14;
  reg signed [32-1:0] _saxi_register_15;
  reg signed [32-1:0] _saxi_register_16;
  reg signed [32-1:0] _saxi_register_17;
  reg signed [32-1:0] _saxi_register_18;
  reg signed [32-1:0] _saxi_register_19;
  reg signed [32-1:0] _saxi_register_20;
  reg signed [32-1:0] _saxi_register_21;
  reg signed [32-1:0] _saxi_register_22;
  reg signed [32-1:0] _saxi_register_23;
  reg signed [32-1:0] _saxi_register_24;
  reg signed [32-1:0] _saxi_register_25;
  reg signed [32-1:0] _saxi_register_26;
  reg signed [32-1:0] _saxi_register_27;
  reg signed [32-1:0] _saxi_register_28;
  reg signed [32-1:0] _saxi_register_29;
  reg signed [32-1:0] _saxi_register_30;
  reg signed [32-1:0] _saxi_register_31;
  reg signed [32-1:0] _saxi_register_32;
  reg signed [32-1:0] _saxi_register_33;
  reg signed [32-1:0] _saxi_register_34;
  reg signed [32-1:0] _saxi_register_35;
  reg signed [32-1:0] _saxi_register_36;
  reg _saxi_flag_0;
  reg _saxi_flag_1;
  reg _saxi_flag_2;
  reg _saxi_flag_3;
  reg _saxi_flag_4;
  reg _saxi_flag_5;
  reg _saxi_flag_6;
  reg _saxi_flag_7;
  reg _saxi_flag_8;
  reg _saxi_flag_9;
  reg _saxi_flag_10;
  reg _saxi_flag_11;
  reg _saxi_flag_12;
  reg _saxi_flag_13;
  reg _saxi_flag_14;
  reg _saxi_flag_15;
  reg _saxi_flag_16;
  reg _saxi_flag_17;
  reg _saxi_flag_18;
  reg _saxi_flag_19;
  reg _saxi_flag_20;
  reg _saxi_flag_21;
  reg _saxi_flag_22;
  reg _saxi_flag_23;
  reg _saxi_flag_24;
  reg _saxi_flag_25;
  reg _saxi_flag_26;
  reg _saxi_flag_27;
  reg _saxi_flag_28;
  reg _saxi_flag_29;
  reg _saxi_flag_30;
  reg _saxi_flag_31;
  reg _saxi_flag_32;
  reg _saxi_flag_33;
  reg _saxi_flag_34;
  reg _saxi_flag_35;
  reg _saxi_flag_36;
  reg signed [32-1:0] _saxi_resetval_0;
  reg signed [32-1:0] _saxi_resetval_1;
  reg signed [32-1:0] _saxi_resetval_2;
  reg signed [32-1:0] _saxi_resetval_3;
  reg signed [32-1:0] _saxi_resetval_4;
  reg signed [32-1:0] _saxi_resetval_5;
  reg signed [32-1:0] _saxi_resetval_6;
  reg signed [32-1:0] _saxi_resetval_7;
  reg signed [32-1:0] _saxi_resetval_8;
  reg signed [32-1:0] _saxi_resetval_9;
  reg signed [32-1:0] _saxi_resetval_10;
  reg signed [32-1:0] _saxi_resetval_11;
  reg signed [32-1:0] _saxi_resetval_12;
  reg signed [32-1:0] _saxi_resetval_13;
  reg signed [32-1:0] _saxi_resetval_14;
  reg signed [32-1:0] _saxi_resetval_15;
  reg signed [32-1:0] _saxi_resetval_16;
  reg signed [32-1:0] _saxi_resetval_17;
  reg signed [32-1:0] _saxi_resetval_18;
  reg signed [32-1:0] _saxi_resetval_19;
  reg signed [32-1:0] _saxi_resetval_20;
  reg signed [32-1:0] _saxi_resetval_21;
  reg signed [32-1:0] _saxi_resetval_22;
  reg signed [32-1:0] _saxi_resetval_23;
  reg signed [32-1:0] _saxi_resetval_24;
  reg signed [32-1:0] _saxi_resetval_25;
  reg signed [32-1:0] _saxi_resetval_26;
  reg signed [32-1:0] _saxi_resetval_27;
  reg signed [32-1:0] _saxi_resetval_28;
  reg signed [32-1:0] _saxi_resetval_29;
  reg signed [32-1:0] _saxi_resetval_30;
  reg signed [32-1:0] _saxi_resetval_31;
  reg signed [32-1:0] _saxi_resetval_32;
  reg signed [32-1:0] _saxi_resetval_33;
  reg signed [32-1:0] _saxi_resetval_34;
  reg signed [32-1:0] _saxi_resetval_35;
  reg signed [32-1:0] _saxi_resetval_36;
  localparam _saxi_maskwidth = 6;
  localparam _saxi_mask = { _saxi_maskwidth{ 1'd1 } };
  localparam _saxi_shift = 2;
  reg [32-1:0] _saxi_register_fsm;
  localparam _saxi_register_fsm_init = 0;
  reg [32-1:0] addr_40;
  reg writevalid_41;
  reg readvalid_42;
  reg prev_awvalid_43;
  reg prev_arvalid_44;
  assign saxi_awready = (_saxi_register_fsm == 0) && (!writevalid_41 && !readvalid_42 && !saxi_bvalid && prev_awvalid_43);
  assign saxi_arready = (_saxi_register_fsm == 0) && (!readvalid_42 && !writevalid_41 && prev_arvalid_44 && !prev_awvalid_43);
  reg [_saxi_maskwidth-1:0] axis_maskaddr_45;
  wire signed [32-1:0] axislite_rdata_46;
  assign axislite_rdata_46 = (axis_maskaddr_45 == 0)? _saxi_register_0 : 
                             (axis_maskaddr_45 == 1)? _saxi_register_1 : 
                             (axis_maskaddr_45 == 2)? _saxi_register_2 : 
                             (axis_maskaddr_45 == 3)? _saxi_register_3 : 
                             (axis_maskaddr_45 == 4)? _saxi_register_4 : 
                             (axis_maskaddr_45 == 5)? _saxi_register_5 : 
                             (axis_maskaddr_45 == 6)? _saxi_register_6 : 
                             (axis_maskaddr_45 == 7)? _saxi_register_7 : 
                             (axis_maskaddr_45 == 8)? _saxi_register_8 : 
                             (axis_maskaddr_45 == 9)? _saxi_register_9 : 
                             (axis_maskaddr_45 == 10)? _saxi_register_10 : 
                             (axis_maskaddr_45 == 11)? _saxi_register_11 : 
                             (axis_maskaddr_45 == 12)? _saxi_register_12 : 
                             (axis_maskaddr_45 == 13)? _saxi_register_13 : 
                             (axis_maskaddr_45 == 14)? _saxi_register_14 : 
                             (axis_maskaddr_45 == 15)? _saxi_register_15 : 
                             (axis_maskaddr_45 == 16)? _saxi_register_16 : 
                             (axis_maskaddr_45 == 17)? _saxi_register_17 : 
                             (axis_maskaddr_45 == 18)? _saxi_register_18 : 
                             (axis_maskaddr_45 == 19)? _saxi_register_19 : 
                             (axis_maskaddr_45 == 20)? _saxi_register_20 : 
                             (axis_maskaddr_45 == 21)? _saxi_register_21 : 
                             (axis_maskaddr_45 == 22)? _saxi_register_22 : 
                             (axis_maskaddr_45 == 23)? _saxi_register_23 : 
                             (axis_maskaddr_45 == 24)? _saxi_register_24 : 
                             (axis_maskaddr_45 == 25)? _saxi_register_25 : 
                             (axis_maskaddr_45 == 26)? _saxi_register_26 : 
                             (axis_maskaddr_45 == 27)? _saxi_register_27 : 
                             (axis_maskaddr_45 == 28)? _saxi_register_28 : 
                             (axis_maskaddr_45 == 29)? _saxi_register_29 : 
                             (axis_maskaddr_45 == 30)? _saxi_register_30 : 
                             (axis_maskaddr_45 == 31)? _saxi_register_31 : 
                             (axis_maskaddr_45 == 32)? _saxi_register_32 : 
                             (axis_maskaddr_45 == 33)? _saxi_register_33 : 
                             (axis_maskaddr_45 == 34)? _saxi_register_34 : 
                             (axis_maskaddr_45 == 35)? _saxi_register_35 : 
                             (axis_maskaddr_45 == 36)? _saxi_register_36 : 'hx;
  wire axislite_flag_47;
  assign axislite_flag_47 = (axis_maskaddr_45 == 0)? _saxi_flag_0 : 
                            (axis_maskaddr_45 == 1)? _saxi_flag_1 : 
                            (axis_maskaddr_45 == 2)? _saxi_flag_2 : 
                            (axis_maskaddr_45 == 3)? _saxi_flag_3 : 
                            (axis_maskaddr_45 == 4)? _saxi_flag_4 : 
                            (axis_maskaddr_45 == 5)? _saxi_flag_5 : 
                            (axis_maskaddr_45 == 6)? _saxi_flag_6 : 
                            (axis_maskaddr_45 == 7)? _saxi_flag_7 : 
                            (axis_maskaddr_45 == 8)? _saxi_flag_8 : 
                            (axis_maskaddr_45 == 9)? _saxi_flag_9 : 
                            (axis_maskaddr_45 == 10)? _saxi_flag_10 : 
                            (axis_maskaddr_45 == 11)? _saxi_flag_11 : 
                            (axis_maskaddr_45 == 12)? _saxi_flag_12 : 
                            (axis_maskaddr_45 == 13)? _saxi_flag_13 : 
                            (axis_maskaddr_45 == 14)? _saxi_flag_14 : 
                            (axis_maskaddr_45 == 15)? _saxi_flag_15 : 
                            (axis_maskaddr_45 == 16)? _saxi_flag_16 : 
                            (axis_maskaddr_45 == 17)? _saxi_flag_17 : 
                            (axis_maskaddr_45 == 18)? _saxi_flag_18 : 
                            (axis_maskaddr_45 == 19)? _saxi_flag_19 : 
                            (axis_maskaddr_45 == 20)? _saxi_flag_20 : 
                            (axis_maskaddr_45 == 21)? _saxi_flag_21 : 
                            (axis_maskaddr_45 == 22)? _saxi_flag_22 : 
                            (axis_maskaddr_45 == 23)? _saxi_flag_23 : 
                            (axis_maskaddr_45 == 24)? _saxi_flag_24 : 
                            (axis_maskaddr_45 == 25)? _saxi_flag_25 : 
                            (axis_maskaddr_45 == 26)? _saxi_flag_26 : 
                            (axis_maskaddr_45 == 27)? _saxi_flag_27 : 
                            (axis_maskaddr_45 == 28)? _saxi_flag_28 : 
                            (axis_maskaddr_45 == 29)? _saxi_flag_29 : 
                            (axis_maskaddr_45 == 30)? _saxi_flag_30 : 
                            (axis_maskaddr_45 == 31)? _saxi_flag_31 : 
                            (axis_maskaddr_45 == 32)? _saxi_flag_32 : 
                            (axis_maskaddr_45 == 33)? _saxi_flag_33 : 
                            (axis_maskaddr_45 == 34)? _saxi_flag_34 : 
                            (axis_maskaddr_45 == 35)? _saxi_flag_35 : 
                            (axis_maskaddr_45 == 36)? _saxi_flag_36 : 'hx;
  wire signed [32-1:0] axislite_resetval_48;
  assign axislite_resetval_48 = (axis_maskaddr_45 == 0)? _saxi_resetval_0 : 
                                (axis_maskaddr_45 == 1)? _saxi_resetval_1 : 
                                (axis_maskaddr_45 == 2)? _saxi_resetval_2 : 
                                (axis_maskaddr_45 == 3)? _saxi_resetval_3 : 
                                (axis_maskaddr_45 == 4)? _saxi_resetval_4 : 
                                (axis_maskaddr_45 == 5)? _saxi_resetval_5 : 
                                (axis_maskaddr_45 == 6)? _saxi_resetval_6 : 
                                (axis_maskaddr_45 == 7)? _saxi_resetval_7 : 
                                (axis_maskaddr_45 == 8)? _saxi_resetval_8 : 
                                (axis_maskaddr_45 == 9)? _saxi_resetval_9 : 
                                (axis_maskaddr_45 == 10)? _saxi_resetval_10 : 
                                (axis_maskaddr_45 == 11)? _saxi_resetval_11 : 
                                (axis_maskaddr_45 == 12)? _saxi_resetval_12 : 
                                (axis_maskaddr_45 == 13)? _saxi_resetval_13 : 
                                (axis_maskaddr_45 == 14)? _saxi_resetval_14 : 
                                (axis_maskaddr_45 == 15)? _saxi_resetval_15 : 
                                (axis_maskaddr_45 == 16)? _saxi_resetval_16 : 
                                (axis_maskaddr_45 == 17)? _saxi_resetval_17 : 
                                (axis_maskaddr_45 == 18)? _saxi_resetval_18 : 
                                (axis_maskaddr_45 == 19)? _saxi_resetval_19 : 
                                (axis_maskaddr_45 == 20)? _saxi_resetval_20 : 
                                (axis_maskaddr_45 == 21)? _saxi_resetval_21 : 
                                (axis_maskaddr_45 == 22)? _saxi_resetval_22 : 
                                (axis_maskaddr_45 == 23)? _saxi_resetval_23 : 
                                (axis_maskaddr_45 == 24)? _saxi_resetval_24 : 
                                (axis_maskaddr_45 == 25)? _saxi_resetval_25 : 
                                (axis_maskaddr_45 == 26)? _saxi_resetval_26 : 
                                (axis_maskaddr_45 == 27)? _saxi_resetval_27 : 
                                (axis_maskaddr_45 == 28)? _saxi_resetval_28 : 
                                (axis_maskaddr_45 == 29)? _saxi_resetval_29 : 
                                (axis_maskaddr_45 == 30)? _saxi_resetval_30 : 
                                (axis_maskaddr_45 == 31)? _saxi_resetval_31 : 
                                (axis_maskaddr_45 == 32)? _saxi_resetval_32 : 
                                (axis_maskaddr_45 == 33)? _saxi_resetval_33 : 
                                (axis_maskaddr_45 == 34)? _saxi_resetval_34 : 
                                (axis_maskaddr_45 == 35)? _saxi_resetval_35 : 
                                (axis_maskaddr_45 == 36)? _saxi_resetval_36 : 'hx;
  reg _saxi_rdata_cond_0_1;
  assign saxi_wready = _saxi_register_fsm == 3;
  wire maxi_idle;
  assign maxi_idle = _maxi_write_idle & _maxi_read_idle;
  wire sw_rst_logic;
  assign sw_rst_logic = maxi_idle & _saxi_register_6;
  wire rst_logic;
  assign rst_logic = RESETN_inv_buf | sw_rst_logic;
  reg RST;
  reg _rst_logic_1;
  reg _rst_logic_2;
  wire signed [32-1:0] irq_49;
  assign irq_49 = _saxi_register_9 & _saxi_register_10;
  wire irq_busy;
  assign irq_busy = _saxi_register_5[0];
  reg irq_busy_edge_50;
  wire irq_busy_edge_51;
  assign irq_busy_edge_51 = irq_busy_edge_50 & !irq_busy;
  wire irq_extern;
  assign irq_extern = |_saxi_register_7;
  reg irq_extern_edge_52;
  wire irq_extern_edge_53;
  assign irq_extern_edge_53 = !irq_extern_edge_52 & irq_extern;
  wire [16-1:0] ram_w8_l262144_id0_0_0_addr;
  wire [8-1:0] ram_w8_l262144_id0_0_0_rdata;
  wire [8-1:0] ram_w8_l262144_id0_0_0_wdata;
  wire ram_w8_l262144_id0_0_0_wenable;
  wire ram_w8_l262144_id0_0_0_enable;
  wire [16-1:0] ram_w8_l262144_id0_0_1_addr;
  wire [8-1:0] ram_w8_l262144_id0_0_1_rdata;
  wire [8-1:0] ram_w8_l262144_id0_0_1_wdata;
  wire ram_w8_l262144_id0_0_1_wenable;
  wire ram_w8_l262144_id0_0_1_enable;
  assign ram_w8_l262144_id0_0_0_wdata = 'hx;
  assign ram_w8_l262144_id0_0_0_wenable = 0;

  ram_w8_l262144_id0_0
  inst_ram_w8_l262144_id0_0
  (
    .CLK(CLK),
    .ram_w8_l262144_id0_0_0_addr(ram_w8_l262144_id0_0_0_addr),
    .ram_w8_l262144_id0_0_0_rdata(ram_w8_l262144_id0_0_0_rdata),
    .ram_w8_l262144_id0_0_0_wdata(ram_w8_l262144_id0_0_0_wdata),
    .ram_w8_l262144_id0_0_0_wenable(ram_w8_l262144_id0_0_0_wenable),
    .ram_w8_l262144_id0_0_0_enable(ram_w8_l262144_id0_0_0_enable),
    .ram_w8_l262144_id0_0_1_addr(ram_w8_l262144_id0_0_1_addr),
    .ram_w8_l262144_id0_0_1_rdata(ram_w8_l262144_id0_0_1_rdata),
    .ram_w8_l262144_id0_0_1_wdata(ram_w8_l262144_id0_0_1_wdata),
    .ram_w8_l262144_id0_0_1_wenable(ram_w8_l262144_id0_0_1_wenable),
    .ram_w8_l262144_id0_0_1_enable(ram_w8_l262144_id0_0_1_enable)
  );

  wire [16-1:0] ram_w8_l262144_id0_1_0_addr;
  wire [8-1:0] ram_w8_l262144_id0_1_0_rdata;
  wire [8-1:0] ram_w8_l262144_id0_1_0_wdata;
  wire ram_w8_l262144_id0_1_0_wenable;
  wire ram_w8_l262144_id0_1_0_enable;
  wire [16-1:0] ram_w8_l262144_id0_1_1_addr;
  wire [8-1:0] ram_w8_l262144_id0_1_1_rdata;
  wire [8-1:0] ram_w8_l262144_id0_1_1_wdata;
  wire ram_w8_l262144_id0_1_1_wenable;
  wire ram_w8_l262144_id0_1_1_enable;
  assign ram_w8_l262144_id0_1_0_wdata = 'hx;
  assign ram_w8_l262144_id0_1_0_wenable = 0;

  ram_w8_l262144_id0_1
  inst_ram_w8_l262144_id0_1
  (
    .CLK(CLK),
    .ram_w8_l262144_id0_1_0_addr(ram_w8_l262144_id0_1_0_addr),
    .ram_w8_l262144_id0_1_0_rdata(ram_w8_l262144_id0_1_0_rdata),
    .ram_w8_l262144_id0_1_0_wdata(ram_w8_l262144_id0_1_0_wdata),
    .ram_w8_l262144_id0_1_0_wenable(ram_w8_l262144_id0_1_0_wenable),
    .ram_w8_l262144_id0_1_0_enable(ram_w8_l262144_id0_1_0_enable),
    .ram_w8_l262144_id0_1_1_addr(ram_w8_l262144_id0_1_1_addr),
    .ram_w8_l262144_id0_1_1_rdata(ram_w8_l262144_id0_1_1_rdata),
    .ram_w8_l262144_id0_1_1_wdata(ram_w8_l262144_id0_1_1_wdata),
    .ram_w8_l262144_id0_1_1_wenable(ram_w8_l262144_id0_1_1_wenable),
    .ram_w8_l262144_id0_1_1_enable(ram_w8_l262144_id0_1_1_enable)
  );

  wire [16-1:0] ram_w8_l262144_id0_2_0_addr;
  wire [8-1:0] ram_w8_l262144_id0_2_0_rdata;
  wire [8-1:0] ram_w8_l262144_id0_2_0_wdata;
  wire ram_w8_l262144_id0_2_0_wenable;
  wire ram_w8_l262144_id0_2_0_enable;
  wire [16-1:0] ram_w8_l262144_id0_2_1_addr;
  wire [8-1:0] ram_w8_l262144_id0_2_1_rdata;
  wire [8-1:0] ram_w8_l262144_id0_2_1_wdata;
  wire ram_w8_l262144_id0_2_1_wenable;
  wire ram_w8_l262144_id0_2_1_enable;
  assign ram_w8_l262144_id0_2_0_wdata = 'hx;
  assign ram_w8_l262144_id0_2_0_wenable = 0;

  ram_w8_l262144_id0_2
  inst_ram_w8_l262144_id0_2
  (
    .CLK(CLK),
    .ram_w8_l262144_id0_2_0_addr(ram_w8_l262144_id0_2_0_addr),
    .ram_w8_l262144_id0_2_0_rdata(ram_w8_l262144_id0_2_0_rdata),
    .ram_w8_l262144_id0_2_0_wdata(ram_w8_l262144_id0_2_0_wdata),
    .ram_w8_l262144_id0_2_0_wenable(ram_w8_l262144_id0_2_0_wenable),
    .ram_w8_l262144_id0_2_0_enable(ram_w8_l262144_id0_2_0_enable),
    .ram_w8_l262144_id0_2_1_addr(ram_w8_l262144_id0_2_1_addr),
    .ram_w8_l262144_id0_2_1_rdata(ram_w8_l262144_id0_2_1_rdata),
    .ram_w8_l262144_id0_2_1_wdata(ram_w8_l262144_id0_2_1_wdata),
    .ram_w8_l262144_id0_2_1_wenable(ram_w8_l262144_id0_2_1_wenable),
    .ram_w8_l262144_id0_2_1_enable(ram_w8_l262144_id0_2_1_enable)
  );

  wire [16-1:0] ram_w8_l262144_id0_3_0_addr;
  wire [8-1:0] ram_w8_l262144_id0_3_0_rdata;
  wire [8-1:0] ram_w8_l262144_id0_3_0_wdata;
  wire ram_w8_l262144_id0_3_0_wenable;
  wire ram_w8_l262144_id0_3_0_enable;
  wire [16-1:0] ram_w8_l262144_id0_3_1_addr;
  wire [8-1:0] ram_w8_l262144_id0_3_1_rdata;
  wire [8-1:0] ram_w8_l262144_id0_3_1_wdata;
  wire ram_w8_l262144_id0_3_1_wenable;
  wire ram_w8_l262144_id0_3_1_enable;
  assign ram_w8_l262144_id0_3_0_wdata = 'hx;
  assign ram_w8_l262144_id0_3_0_wenable = 0;

  ram_w8_l262144_id0_3
  inst_ram_w8_l262144_id0_3
  (
    .CLK(CLK),
    .ram_w8_l262144_id0_3_0_addr(ram_w8_l262144_id0_3_0_addr),
    .ram_w8_l262144_id0_3_0_rdata(ram_w8_l262144_id0_3_0_rdata),
    .ram_w8_l262144_id0_3_0_wdata(ram_w8_l262144_id0_3_0_wdata),
    .ram_w8_l262144_id0_3_0_wenable(ram_w8_l262144_id0_3_0_wenable),
    .ram_w8_l262144_id0_3_0_enable(ram_w8_l262144_id0_3_0_enable),
    .ram_w8_l262144_id0_3_1_addr(ram_w8_l262144_id0_3_1_addr),
    .ram_w8_l262144_id0_3_1_rdata(ram_w8_l262144_id0_3_1_rdata),
    .ram_w8_l262144_id0_3_1_wdata(ram_w8_l262144_id0_3_1_wdata),
    .ram_w8_l262144_id0_3_1_wenable(ram_w8_l262144_id0_3_1_wenable),
    .ram_w8_l262144_id0_3_1_enable(ram_w8_l262144_id0_3_1_enable)
  );

  wire [13-1:0] ram_w8_l32768_id0_0_0_addr;
  wire [8-1:0] ram_w8_l32768_id0_0_0_rdata;
  wire [8-1:0] ram_w8_l32768_id0_0_0_wdata;
  wire ram_w8_l32768_id0_0_0_wenable;
  wire ram_w8_l32768_id0_0_0_enable;
  wire [13-1:0] ram_w8_l32768_id0_0_1_addr;
  wire [8-1:0] ram_w8_l32768_id0_0_1_rdata;
  wire [8-1:0] ram_w8_l32768_id0_0_1_wdata;
  wire ram_w8_l32768_id0_0_1_wenable;
  wire ram_w8_l32768_id0_0_1_enable;
  assign ram_w8_l32768_id0_0_0_wdata = 'hx;
  assign ram_w8_l32768_id0_0_0_wenable = 0;

  ram_w8_l32768_id0_0
  inst_ram_w8_l32768_id0_0
  (
    .CLK(CLK),
    .ram_w8_l32768_id0_0_0_addr(ram_w8_l32768_id0_0_0_addr),
    .ram_w8_l32768_id0_0_0_rdata(ram_w8_l32768_id0_0_0_rdata),
    .ram_w8_l32768_id0_0_0_wdata(ram_w8_l32768_id0_0_0_wdata),
    .ram_w8_l32768_id0_0_0_wenable(ram_w8_l32768_id0_0_0_wenable),
    .ram_w8_l32768_id0_0_0_enable(ram_w8_l32768_id0_0_0_enable),
    .ram_w8_l32768_id0_0_1_addr(ram_w8_l32768_id0_0_1_addr),
    .ram_w8_l32768_id0_0_1_rdata(ram_w8_l32768_id0_0_1_rdata),
    .ram_w8_l32768_id0_0_1_wdata(ram_w8_l32768_id0_0_1_wdata),
    .ram_w8_l32768_id0_0_1_wenable(ram_w8_l32768_id0_0_1_wenable),
    .ram_w8_l32768_id0_0_1_enable(ram_w8_l32768_id0_0_1_enable)
  );

  wire [13-1:0] ram_w8_l32768_id0_1_0_addr;
  wire [8-1:0] ram_w8_l32768_id0_1_0_rdata;
  wire [8-1:0] ram_w8_l32768_id0_1_0_wdata;
  wire ram_w8_l32768_id0_1_0_wenable;
  wire ram_w8_l32768_id0_1_0_enable;
  wire [13-1:0] ram_w8_l32768_id0_1_1_addr;
  wire [8-1:0] ram_w8_l32768_id0_1_1_rdata;
  wire [8-1:0] ram_w8_l32768_id0_1_1_wdata;
  wire ram_w8_l32768_id0_1_1_wenable;
  wire ram_w8_l32768_id0_1_1_enable;
  assign ram_w8_l32768_id0_1_0_wdata = 'hx;
  assign ram_w8_l32768_id0_1_0_wenable = 0;

  ram_w8_l32768_id0_1
  inst_ram_w8_l32768_id0_1
  (
    .CLK(CLK),
    .ram_w8_l32768_id0_1_0_addr(ram_w8_l32768_id0_1_0_addr),
    .ram_w8_l32768_id0_1_0_rdata(ram_w8_l32768_id0_1_0_rdata),
    .ram_w8_l32768_id0_1_0_wdata(ram_w8_l32768_id0_1_0_wdata),
    .ram_w8_l32768_id0_1_0_wenable(ram_w8_l32768_id0_1_0_wenable),
    .ram_w8_l32768_id0_1_0_enable(ram_w8_l32768_id0_1_0_enable),
    .ram_w8_l32768_id0_1_1_addr(ram_w8_l32768_id0_1_1_addr),
    .ram_w8_l32768_id0_1_1_rdata(ram_w8_l32768_id0_1_1_rdata),
    .ram_w8_l32768_id0_1_1_wdata(ram_w8_l32768_id0_1_1_wdata),
    .ram_w8_l32768_id0_1_1_wenable(ram_w8_l32768_id0_1_1_wenable),
    .ram_w8_l32768_id0_1_1_enable(ram_w8_l32768_id0_1_1_enable)
  );

  wire [13-1:0] ram_w8_l32768_id0_2_0_addr;
  wire [8-1:0] ram_w8_l32768_id0_2_0_rdata;
  wire [8-1:0] ram_w8_l32768_id0_2_0_wdata;
  wire ram_w8_l32768_id0_2_0_wenable;
  wire ram_w8_l32768_id0_2_0_enable;
  wire [13-1:0] ram_w8_l32768_id0_2_1_addr;
  wire [8-1:0] ram_w8_l32768_id0_2_1_rdata;
  wire [8-1:0] ram_w8_l32768_id0_2_1_wdata;
  wire ram_w8_l32768_id0_2_1_wenable;
  wire ram_w8_l32768_id0_2_1_enable;
  assign ram_w8_l32768_id0_2_0_wdata = 'hx;
  assign ram_w8_l32768_id0_2_0_wenable = 0;

  ram_w8_l32768_id0_2
  inst_ram_w8_l32768_id0_2
  (
    .CLK(CLK),
    .ram_w8_l32768_id0_2_0_addr(ram_w8_l32768_id0_2_0_addr),
    .ram_w8_l32768_id0_2_0_rdata(ram_w8_l32768_id0_2_0_rdata),
    .ram_w8_l32768_id0_2_0_wdata(ram_w8_l32768_id0_2_0_wdata),
    .ram_w8_l32768_id0_2_0_wenable(ram_w8_l32768_id0_2_0_wenable),
    .ram_w8_l32768_id0_2_0_enable(ram_w8_l32768_id0_2_0_enable),
    .ram_w8_l32768_id0_2_1_addr(ram_w8_l32768_id0_2_1_addr),
    .ram_w8_l32768_id0_2_1_rdata(ram_w8_l32768_id0_2_1_rdata),
    .ram_w8_l32768_id0_2_1_wdata(ram_w8_l32768_id0_2_1_wdata),
    .ram_w8_l32768_id0_2_1_wenable(ram_w8_l32768_id0_2_1_wenable),
    .ram_w8_l32768_id0_2_1_enable(ram_w8_l32768_id0_2_1_enable)
  );

  wire [13-1:0] ram_w8_l32768_id0_3_0_addr;
  wire [8-1:0] ram_w8_l32768_id0_3_0_rdata;
  wire [8-1:0] ram_w8_l32768_id0_3_0_wdata;
  wire ram_w8_l32768_id0_3_0_wenable;
  wire ram_w8_l32768_id0_3_0_enable;
  wire [13-1:0] ram_w8_l32768_id0_3_1_addr;
  wire [8-1:0] ram_w8_l32768_id0_3_1_rdata;
  wire [8-1:0] ram_w8_l32768_id0_3_1_wdata;
  wire ram_w8_l32768_id0_3_1_wenable;
  wire ram_w8_l32768_id0_3_1_enable;
  assign ram_w8_l32768_id0_3_0_wdata = 'hx;
  assign ram_w8_l32768_id0_3_0_wenable = 0;

  ram_w8_l32768_id0_3
  inst_ram_w8_l32768_id0_3
  (
    .CLK(CLK),
    .ram_w8_l32768_id0_3_0_addr(ram_w8_l32768_id0_3_0_addr),
    .ram_w8_l32768_id0_3_0_rdata(ram_w8_l32768_id0_3_0_rdata),
    .ram_w8_l32768_id0_3_0_wdata(ram_w8_l32768_id0_3_0_wdata),
    .ram_w8_l32768_id0_3_0_wenable(ram_w8_l32768_id0_3_0_wenable),
    .ram_w8_l32768_id0_3_0_enable(ram_w8_l32768_id0_3_0_enable),
    .ram_w8_l32768_id0_3_1_addr(ram_w8_l32768_id0_3_1_addr),
    .ram_w8_l32768_id0_3_1_rdata(ram_w8_l32768_id0_3_1_rdata),
    .ram_w8_l32768_id0_3_1_wdata(ram_w8_l32768_id0_3_1_wdata),
    .ram_w8_l32768_id0_3_1_wenable(ram_w8_l32768_id0_3_1_wenable),
    .ram_w8_l32768_id0_3_1_enable(ram_w8_l32768_id0_3_1_enable)
  );

  wire [12-1:0] ram_w8_l16384_id0_0_0_addr;
  wire [8-1:0] ram_w8_l16384_id0_0_0_rdata;
  wire [8-1:0] ram_w8_l16384_id0_0_0_wdata;
  wire ram_w8_l16384_id0_0_0_wenable;
  wire ram_w8_l16384_id0_0_0_enable;
  wire [12-1:0] ram_w8_l16384_id0_0_1_addr;
  wire [8-1:0] ram_w8_l16384_id0_0_1_rdata;
  wire [8-1:0] ram_w8_l16384_id0_0_1_wdata;
  wire ram_w8_l16384_id0_0_1_wenable;
  wire ram_w8_l16384_id0_0_1_enable;

  ram_w8_l16384_id0_0
  inst_ram_w8_l16384_id0_0
  (
    .CLK(CLK),
    .ram_w8_l16384_id0_0_0_addr(ram_w8_l16384_id0_0_0_addr),
    .ram_w8_l16384_id0_0_0_rdata(ram_w8_l16384_id0_0_0_rdata),
    .ram_w8_l16384_id0_0_0_wdata(ram_w8_l16384_id0_0_0_wdata),
    .ram_w8_l16384_id0_0_0_wenable(ram_w8_l16384_id0_0_0_wenable),
    .ram_w8_l16384_id0_0_0_enable(ram_w8_l16384_id0_0_0_enable),
    .ram_w8_l16384_id0_0_1_addr(ram_w8_l16384_id0_0_1_addr),
    .ram_w8_l16384_id0_0_1_rdata(ram_w8_l16384_id0_0_1_rdata),
    .ram_w8_l16384_id0_0_1_wdata(ram_w8_l16384_id0_0_1_wdata),
    .ram_w8_l16384_id0_0_1_wenable(ram_w8_l16384_id0_0_1_wenable),
    .ram_w8_l16384_id0_0_1_enable(ram_w8_l16384_id0_0_1_enable)
  );

  wire [12-1:0] ram_w8_l16384_id0_1_0_addr;
  wire [8-1:0] ram_w8_l16384_id0_1_0_rdata;
  wire [8-1:0] ram_w8_l16384_id0_1_0_wdata;
  wire ram_w8_l16384_id0_1_0_wenable;
  wire ram_w8_l16384_id0_1_0_enable;
  wire [12-1:0] ram_w8_l16384_id0_1_1_addr;
  wire [8-1:0] ram_w8_l16384_id0_1_1_rdata;
  wire [8-1:0] ram_w8_l16384_id0_1_1_wdata;
  wire ram_w8_l16384_id0_1_1_wenable;
  wire ram_w8_l16384_id0_1_1_enable;

  ram_w8_l16384_id0_1
  inst_ram_w8_l16384_id0_1
  (
    .CLK(CLK),
    .ram_w8_l16384_id0_1_0_addr(ram_w8_l16384_id0_1_0_addr),
    .ram_w8_l16384_id0_1_0_rdata(ram_w8_l16384_id0_1_0_rdata),
    .ram_w8_l16384_id0_1_0_wdata(ram_w8_l16384_id0_1_0_wdata),
    .ram_w8_l16384_id0_1_0_wenable(ram_w8_l16384_id0_1_0_wenable),
    .ram_w8_l16384_id0_1_0_enable(ram_w8_l16384_id0_1_0_enable),
    .ram_w8_l16384_id0_1_1_addr(ram_w8_l16384_id0_1_1_addr),
    .ram_w8_l16384_id0_1_1_rdata(ram_w8_l16384_id0_1_1_rdata),
    .ram_w8_l16384_id0_1_1_wdata(ram_w8_l16384_id0_1_1_wdata),
    .ram_w8_l16384_id0_1_1_wenable(ram_w8_l16384_id0_1_1_wenable),
    .ram_w8_l16384_id0_1_1_enable(ram_w8_l16384_id0_1_1_enable)
  );

  wire [12-1:0] ram_w8_l16384_id0_2_0_addr;
  wire [8-1:0] ram_w8_l16384_id0_2_0_rdata;
  wire [8-1:0] ram_w8_l16384_id0_2_0_wdata;
  wire ram_w8_l16384_id0_2_0_wenable;
  wire ram_w8_l16384_id0_2_0_enable;
  wire [12-1:0] ram_w8_l16384_id0_2_1_addr;
  wire [8-1:0] ram_w8_l16384_id0_2_1_rdata;
  wire [8-1:0] ram_w8_l16384_id0_2_1_wdata;
  wire ram_w8_l16384_id0_2_1_wenable;
  wire ram_w8_l16384_id0_2_1_enable;

  ram_w8_l16384_id0_2
  inst_ram_w8_l16384_id0_2
  (
    .CLK(CLK),
    .ram_w8_l16384_id0_2_0_addr(ram_w8_l16384_id0_2_0_addr),
    .ram_w8_l16384_id0_2_0_rdata(ram_w8_l16384_id0_2_0_rdata),
    .ram_w8_l16384_id0_2_0_wdata(ram_w8_l16384_id0_2_0_wdata),
    .ram_w8_l16384_id0_2_0_wenable(ram_w8_l16384_id0_2_0_wenable),
    .ram_w8_l16384_id0_2_0_enable(ram_w8_l16384_id0_2_0_enable),
    .ram_w8_l16384_id0_2_1_addr(ram_w8_l16384_id0_2_1_addr),
    .ram_w8_l16384_id0_2_1_rdata(ram_w8_l16384_id0_2_1_rdata),
    .ram_w8_l16384_id0_2_1_wdata(ram_w8_l16384_id0_2_1_wdata),
    .ram_w8_l16384_id0_2_1_wenable(ram_w8_l16384_id0_2_1_wenable),
    .ram_w8_l16384_id0_2_1_enable(ram_w8_l16384_id0_2_1_enable)
  );

  wire [12-1:0] ram_w8_l16384_id0_3_0_addr;
  wire [8-1:0] ram_w8_l16384_id0_3_0_rdata;
  wire [8-1:0] ram_w8_l16384_id0_3_0_wdata;
  wire ram_w8_l16384_id0_3_0_wenable;
  wire ram_w8_l16384_id0_3_0_enable;
  wire [12-1:0] ram_w8_l16384_id0_3_1_addr;
  wire [8-1:0] ram_w8_l16384_id0_3_1_rdata;
  wire [8-1:0] ram_w8_l16384_id0_3_1_wdata;
  wire ram_w8_l16384_id0_3_1_wenable;
  wire ram_w8_l16384_id0_3_1_enable;

  ram_w8_l16384_id0_3
  inst_ram_w8_l16384_id0_3
  (
    .CLK(CLK),
    .ram_w8_l16384_id0_3_0_addr(ram_w8_l16384_id0_3_0_addr),
    .ram_w8_l16384_id0_3_0_rdata(ram_w8_l16384_id0_3_0_rdata),
    .ram_w8_l16384_id0_3_0_wdata(ram_w8_l16384_id0_3_0_wdata),
    .ram_w8_l16384_id0_3_0_wenable(ram_w8_l16384_id0_3_0_wenable),
    .ram_w8_l16384_id0_3_0_enable(ram_w8_l16384_id0_3_0_enable),
    .ram_w8_l16384_id0_3_1_addr(ram_w8_l16384_id0_3_1_addr),
    .ram_w8_l16384_id0_3_1_rdata(ram_w8_l16384_id0_3_1_rdata),
    .ram_w8_l16384_id0_3_1_wdata(ram_w8_l16384_id0_3_1_wdata),
    .ram_w8_l16384_id0_3_1_wenable(ram_w8_l16384_id0_3_1_wenable),
    .ram_w8_l16384_id0_3_1_enable(ram_w8_l16384_id0_3_1_enable)
  );

  wire [12-1:0] ram_w8_l16384_id1_0_0_addr;
  wire [8-1:0] ram_w8_l16384_id1_0_0_rdata;
  wire [8-1:0] ram_w8_l16384_id1_0_0_wdata;
  wire ram_w8_l16384_id1_0_0_wenable;
  wire ram_w8_l16384_id1_0_0_enable;
  wire [12-1:0] ram_w8_l16384_id1_0_1_addr;
  wire [8-1:0] ram_w8_l16384_id1_0_1_rdata;
  wire [8-1:0] ram_w8_l16384_id1_0_1_wdata;
  wire ram_w8_l16384_id1_0_1_wenable;
  wire ram_w8_l16384_id1_0_1_enable;

  ram_w8_l16384_id1_0
  inst_ram_w8_l16384_id1_0
  (
    .CLK(CLK),
    .ram_w8_l16384_id1_0_0_addr(ram_w8_l16384_id1_0_0_addr),
    .ram_w8_l16384_id1_0_0_rdata(ram_w8_l16384_id1_0_0_rdata),
    .ram_w8_l16384_id1_0_0_wdata(ram_w8_l16384_id1_0_0_wdata),
    .ram_w8_l16384_id1_0_0_wenable(ram_w8_l16384_id1_0_0_wenable),
    .ram_w8_l16384_id1_0_0_enable(ram_w8_l16384_id1_0_0_enable),
    .ram_w8_l16384_id1_0_1_addr(ram_w8_l16384_id1_0_1_addr),
    .ram_w8_l16384_id1_0_1_rdata(ram_w8_l16384_id1_0_1_rdata),
    .ram_w8_l16384_id1_0_1_wdata(ram_w8_l16384_id1_0_1_wdata),
    .ram_w8_l16384_id1_0_1_wenable(ram_w8_l16384_id1_0_1_wenable),
    .ram_w8_l16384_id1_0_1_enable(ram_w8_l16384_id1_0_1_enable)
  );

  wire [12-1:0] ram_w8_l16384_id1_1_0_addr;
  wire [8-1:0] ram_w8_l16384_id1_1_0_rdata;
  wire [8-1:0] ram_w8_l16384_id1_1_0_wdata;
  wire ram_w8_l16384_id1_1_0_wenable;
  wire ram_w8_l16384_id1_1_0_enable;
  wire [12-1:0] ram_w8_l16384_id1_1_1_addr;
  wire [8-1:0] ram_w8_l16384_id1_1_1_rdata;
  wire [8-1:0] ram_w8_l16384_id1_1_1_wdata;
  wire ram_w8_l16384_id1_1_1_wenable;
  wire ram_w8_l16384_id1_1_1_enable;

  ram_w8_l16384_id1_1
  inst_ram_w8_l16384_id1_1
  (
    .CLK(CLK),
    .ram_w8_l16384_id1_1_0_addr(ram_w8_l16384_id1_1_0_addr),
    .ram_w8_l16384_id1_1_0_rdata(ram_w8_l16384_id1_1_0_rdata),
    .ram_w8_l16384_id1_1_0_wdata(ram_w8_l16384_id1_1_0_wdata),
    .ram_w8_l16384_id1_1_0_wenable(ram_w8_l16384_id1_1_0_wenable),
    .ram_w8_l16384_id1_1_0_enable(ram_w8_l16384_id1_1_0_enable),
    .ram_w8_l16384_id1_1_1_addr(ram_w8_l16384_id1_1_1_addr),
    .ram_w8_l16384_id1_1_1_rdata(ram_w8_l16384_id1_1_1_rdata),
    .ram_w8_l16384_id1_1_1_wdata(ram_w8_l16384_id1_1_1_wdata),
    .ram_w8_l16384_id1_1_1_wenable(ram_w8_l16384_id1_1_1_wenable),
    .ram_w8_l16384_id1_1_1_enable(ram_w8_l16384_id1_1_1_enable)
  );

  wire [12-1:0] ram_w8_l16384_id1_2_0_addr;
  wire [8-1:0] ram_w8_l16384_id1_2_0_rdata;
  wire [8-1:0] ram_w8_l16384_id1_2_0_wdata;
  wire ram_w8_l16384_id1_2_0_wenable;
  wire ram_w8_l16384_id1_2_0_enable;
  wire [12-1:0] ram_w8_l16384_id1_2_1_addr;
  wire [8-1:0] ram_w8_l16384_id1_2_1_rdata;
  wire [8-1:0] ram_w8_l16384_id1_2_1_wdata;
  wire ram_w8_l16384_id1_2_1_wenable;
  wire ram_w8_l16384_id1_2_1_enable;

  ram_w8_l16384_id1_2
  inst_ram_w8_l16384_id1_2
  (
    .CLK(CLK),
    .ram_w8_l16384_id1_2_0_addr(ram_w8_l16384_id1_2_0_addr),
    .ram_w8_l16384_id1_2_0_rdata(ram_w8_l16384_id1_2_0_rdata),
    .ram_w8_l16384_id1_2_0_wdata(ram_w8_l16384_id1_2_0_wdata),
    .ram_w8_l16384_id1_2_0_wenable(ram_w8_l16384_id1_2_0_wenable),
    .ram_w8_l16384_id1_2_0_enable(ram_w8_l16384_id1_2_0_enable),
    .ram_w8_l16384_id1_2_1_addr(ram_w8_l16384_id1_2_1_addr),
    .ram_w8_l16384_id1_2_1_rdata(ram_w8_l16384_id1_2_1_rdata),
    .ram_w8_l16384_id1_2_1_wdata(ram_w8_l16384_id1_2_1_wdata),
    .ram_w8_l16384_id1_2_1_wenable(ram_w8_l16384_id1_2_1_wenable),
    .ram_w8_l16384_id1_2_1_enable(ram_w8_l16384_id1_2_1_enable)
  );

  wire [12-1:0] ram_w8_l16384_id1_3_0_addr;
  wire [8-1:0] ram_w8_l16384_id1_3_0_rdata;
  wire [8-1:0] ram_w8_l16384_id1_3_0_wdata;
  wire ram_w8_l16384_id1_3_0_wenable;
  wire ram_w8_l16384_id1_3_0_enable;
  wire [12-1:0] ram_w8_l16384_id1_3_1_addr;
  wire [8-1:0] ram_w8_l16384_id1_3_1_rdata;
  wire [8-1:0] ram_w8_l16384_id1_3_1_wdata;
  wire ram_w8_l16384_id1_3_1_wenable;
  wire ram_w8_l16384_id1_3_1_enable;

  ram_w8_l16384_id1_3
  inst_ram_w8_l16384_id1_3
  (
    .CLK(CLK),
    .ram_w8_l16384_id1_3_0_addr(ram_w8_l16384_id1_3_0_addr),
    .ram_w8_l16384_id1_3_0_rdata(ram_w8_l16384_id1_3_0_rdata),
    .ram_w8_l16384_id1_3_0_wdata(ram_w8_l16384_id1_3_0_wdata),
    .ram_w8_l16384_id1_3_0_wenable(ram_w8_l16384_id1_3_0_wenable),
    .ram_w8_l16384_id1_3_0_enable(ram_w8_l16384_id1_3_0_enable),
    .ram_w8_l16384_id1_3_1_addr(ram_w8_l16384_id1_3_1_addr),
    .ram_w8_l16384_id1_3_1_rdata(ram_w8_l16384_id1_3_1_rdata),
    .ram_w8_l16384_id1_3_1_wdata(ram_w8_l16384_id1_3_1_wdata),
    .ram_w8_l16384_id1_3_1_wenable(ram_w8_l16384_id1_3_1_wenable),
    .ram_w8_l16384_id1_3_1_enable(ram_w8_l16384_id1_3_1_enable)
  );

  wire [12-1:0] ram_w8_l16384_id2_0_0_addr;
  wire [8-1:0] ram_w8_l16384_id2_0_0_rdata;
  wire [8-1:0] ram_w8_l16384_id2_0_0_wdata;
  wire ram_w8_l16384_id2_0_0_wenable;
  wire ram_w8_l16384_id2_0_0_enable;
  wire [12-1:0] ram_w8_l16384_id2_0_1_addr;
  wire [8-1:0] ram_w8_l16384_id2_0_1_rdata;
  wire [8-1:0] ram_w8_l16384_id2_0_1_wdata;
  wire ram_w8_l16384_id2_0_1_wenable;
  wire ram_w8_l16384_id2_0_1_enable;
  assign ram_w8_l16384_id2_0_0_wdata = 'hx;
  assign ram_w8_l16384_id2_0_0_wenable = 0;

  ram_w8_l16384_id2_0
  inst_ram_w8_l16384_id2_0
  (
    .CLK(CLK),
    .ram_w8_l16384_id2_0_0_addr(ram_w8_l16384_id2_0_0_addr),
    .ram_w8_l16384_id2_0_0_rdata(ram_w8_l16384_id2_0_0_rdata),
    .ram_w8_l16384_id2_0_0_wdata(ram_w8_l16384_id2_0_0_wdata),
    .ram_w8_l16384_id2_0_0_wenable(ram_w8_l16384_id2_0_0_wenable),
    .ram_w8_l16384_id2_0_0_enable(ram_w8_l16384_id2_0_0_enable),
    .ram_w8_l16384_id2_0_1_addr(ram_w8_l16384_id2_0_1_addr),
    .ram_w8_l16384_id2_0_1_rdata(ram_w8_l16384_id2_0_1_rdata),
    .ram_w8_l16384_id2_0_1_wdata(ram_w8_l16384_id2_0_1_wdata),
    .ram_w8_l16384_id2_0_1_wenable(ram_w8_l16384_id2_0_1_wenable),
    .ram_w8_l16384_id2_0_1_enable(ram_w8_l16384_id2_0_1_enable)
  );

  wire [12-1:0] ram_w8_l16384_id2_1_0_addr;
  wire [8-1:0] ram_w8_l16384_id2_1_0_rdata;
  wire [8-1:0] ram_w8_l16384_id2_1_0_wdata;
  wire ram_w8_l16384_id2_1_0_wenable;
  wire ram_w8_l16384_id2_1_0_enable;
  wire [12-1:0] ram_w8_l16384_id2_1_1_addr;
  wire [8-1:0] ram_w8_l16384_id2_1_1_rdata;
  wire [8-1:0] ram_w8_l16384_id2_1_1_wdata;
  wire ram_w8_l16384_id2_1_1_wenable;
  wire ram_w8_l16384_id2_1_1_enable;
  assign ram_w8_l16384_id2_1_0_wdata = 'hx;
  assign ram_w8_l16384_id2_1_0_wenable = 0;

  ram_w8_l16384_id2_1
  inst_ram_w8_l16384_id2_1
  (
    .CLK(CLK),
    .ram_w8_l16384_id2_1_0_addr(ram_w8_l16384_id2_1_0_addr),
    .ram_w8_l16384_id2_1_0_rdata(ram_w8_l16384_id2_1_0_rdata),
    .ram_w8_l16384_id2_1_0_wdata(ram_w8_l16384_id2_1_0_wdata),
    .ram_w8_l16384_id2_1_0_wenable(ram_w8_l16384_id2_1_0_wenable),
    .ram_w8_l16384_id2_1_0_enable(ram_w8_l16384_id2_1_0_enable),
    .ram_w8_l16384_id2_1_1_addr(ram_w8_l16384_id2_1_1_addr),
    .ram_w8_l16384_id2_1_1_rdata(ram_w8_l16384_id2_1_1_rdata),
    .ram_w8_l16384_id2_1_1_wdata(ram_w8_l16384_id2_1_1_wdata),
    .ram_w8_l16384_id2_1_1_wenable(ram_w8_l16384_id2_1_1_wenable),
    .ram_w8_l16384_id2_1_1_enable(ram_w8_l16384_id2_1_1_enable)
  );

  wire [12-1:0] ram_w8_l16384_id2_2_0_addr;
  wire [8-1:0] ram_w8_l16384_id2_2_0_rdata;
  wire [8-1:0] ram_w8_l16384_id2_2_0_wdata;
  wire ram_w8_l16384_id2_2_0_wenable;
  wire ram_w8_l16384_id2_2_0_enable;
  wire [12-1:0] ram_w8_l16384_id2_2_1_addr;
  wire [8-1:0] ram_w8_l16384_id2_2_1_rdata;
  wire [8-1:0] ram_w8_l16384_id2_2_1_wdata;
  wire ram_w8_l16384_id2_2_1_wenable;
  wire ram_w8_l16384_id2_2_1_enable;
  assign ram_w8_l16384_id2_2_0_wdata = 'hx;
  assign ram_w8_l16384_id2_2_0_wenable = 0;

  ram_w8_l16384_id2_2
  inst_ram_w8_l16384_id2_2
  (
    .CLK(CLK),
    .ram_w8_l16384_id2_2_0_addr(ram_w8_l16384_id2_2_0_addr),
    .ram_w8_l16384_id2_2_0_rdata(ram_w8_l16384_id2_2_0_rdata),
    .ram_w8_l16384_id2_2_0_wdata(ram_w8_l16384_id2_2_0_wdata),
    .ram_w8_l16384_id2_2_0_wenable(ram_w8_l16384_id2_2_0_wenable),
    .ram_w8_l16384_id2_2_0_enable(ram_w8_l16384_id2_2_0_enable),
    .ram_w8_l16384_id2_2_1_addr(ram_w8_l16384_id2_2_1_addr),
    .ram_w8_l16384_id2_2_1_rdata(ram_w8_l16384_id2_2_1_rdata),
    .ram_w8_l16384_id2_2_1_wdata(ram_w8_l16384_id2_2_1_wdata),
    .ram_w8_l16384_id2_2_1_wenable(ram_w8_l16384_id2_2_1_wenable),
    .ram_w8_l16384_id2_2_1_enable(ram_w8_l16384_id2_2_1_enable)
  );

  wire [12-1:0] ram_w8_l16384_id2_3_0_addr;
  wire [8-1:0] ram_w8_l16384_id2_3_0_rdata;
  wire [8-1:0] ram_w8_l16384_id2_3_0_wdata;
  wire ram_w8_l16384_id2_3_0_wenable;
  wire ram_w8_l16384_id2_3_0_enable;
  wire [12-1:0] ram_w8_l16384_id2_3_1_addr;
  wire [8-1:0] ram_w8_l16384_id2_3_1_rdata;
  wire [8-1:0] ram_w8_l16384_id2_3_1_wdata;
  wire ram_w8_l16384_id2_3_1_wenable;
  wire ram_w8_l16384_id2_3_1_enable;
  assign ram_w8_l16384_id2_3_0_wdata = 'hx;
  assign ram_w8_l16384_id2_3_0_wenable = 0;

  ram_w8_l16384_id2_3
  inst_ram_w8_l16384_id2_3
  (
    .CLK(CLK),
    .ram_w8_l16384_id2_3_0_addr(ram_w8_l16384_id2_3_0_addr),
    .ram_w8_l16384_id2_3_0_rdata(ram_w8_l16384_id2_3_0_rdata),
    .ram_w8_l16384_id2_3_0_wdata(ram_w8_l16384_id2_3_0_wdata),
    .ram_w8_l16384_id2_3_0_wenable(ram_w8_l16384_id2_3_0_wenable),
    .ram_w8_l16384_id2_3_0_enable(ram_w8_l16384_id2_3_0_enable),
    .ram_w8_l16384_id2_3_1_addr(ram_w8_l16384_id2_3_1_addr),
    .ram_w8_l16384_id2_3_1_rdata(ram_w8_l16384_id2_3_1_rdata),
    .ram_w8_l16384_id2_3_1_wdata(ram_w8_l16384_id2_3_1_wdata),
    .ram_w8_l16384_id2_3_1_wenable(ram_w8_l16384_id2_3_1_wenable),
    .ram_w8_l16384_id2_3_1_enable(ram_w8_l16384_id2_3_1_enable)
  );

  wire [12-1:0] ram_w8_l16384_id3_0_0_addr;
  wire [8-1:0] ram_w8_l16384_id3_0_0_rdata;
  wire [8-1:0] ram_w8_l16384_id3_0_0_wdata;
  wire ram_w8_l16384_id3_0_0_wenable;
  wire ram_w8_l16384_id3_0_0_enable;
  wire [12-1:0] ram_w8_l16384_id3_0_1_addr;
  wire [8-1:0] ram_w8_l16384_id3_0_1_rdata;
  wire [8-1:0] ram_w8_l16384_id3_0_1_wdata;
  wire ram_w8_l16384_id3_0_1_wenable;
  wire ram_w8_l16384_id3_0_1_enable;
  assign ram_w8_l16384_id3_0_0_wdata = 'hx;
  assign ram_w8_l16384_id3_0_0_wenable = 0;

  ram_w8_l16384_id3_0
  inst_ram_w8_l16384_id3_0
  (
    .CLK(CLK),
    .ram_w8_l16384_id3_0_0_addr(ram_w8_l16384_id3_0_0_addr),
    .ram_w8_l16384_id3_0_0_rdata(ram_w8_l16384_id3_0_0_rdata),
    .ram_w8_l16384_id3_0_0_wdata(ram_w8_l16384_id3_0_0_wdata),
    .ram_w8_l16384_id3_0_0_wenable(ram_w8_l16384_id3_0_0_wenable),
    .ram_w8_l16384_id3_0_0_enable(ram_w8_l16384_id3_0_0_enable),
    .ram_w8_l16384_id3_0_1_addr(ram_w8_l16384_id3_0_1_addr),
    .ram_w8_l16384_id3_0_1_rdata(ram_w8_l16384_id3_0_1_rdata),
    .ram_w8_l16384_id3_0_1_wdata(ram_w8_l16384_id3_0_1_wdata),
    .ram_w8_l16384_id3_0_1_wenable(ram_w8_l16384_id3_0_1_wenable),
    .ram_w8_l16384_id3_0_1_enable(ram_w8_l16384_id3_0_1_enable)
  );

  wire [12-1:0] ram_w8_l16384_id3_1_0_addr;
  wire [8-1:0] ram_w8_l16384_id3_1_0_rdata;
  wire [8-1:0] ram_w8_l16384_id3_1_0_wdata;
  wire ram_w8_l16384_id3_1_0_wenable;
  wire ram_w8_l16384_id3_1_0_enable;
  wire [12-1:0] ram_w8_l16384_id3_1_1_addr;
  wire [8-1:0] ram_w8_l16384_id3_1_1_rdata;
  wire [8-1:0] ram_w8_l16384_id3_1_1_wdata;
  wire ram_w8_l16384_id3_1_1_wenable;
  wire ram_w8_l16384_id3_1_1_enable;
  assign ram_w8_l16384_id3_1_0_wdata = 'hx;
  assign ram_w8_l16384_id3_1_0_wenable = 0;

  ram_w8_l16384_id3_1
  inst_ram_w8_l16384_id3_1
  (
    .CLK(CLK),
    .ram_w8_l16384_id3_1_0_addr(ram_w8_l16384_id3_1_0_addr),
    .ram_w8_l16384_id3_1_0_rdata(ram_w8_l16384_id3_1_0_rdata),
    .ram_w8_l16384_id3_1_0_wdata(ram_w8_l16384_id3_1_0_wdata),
    .ram_w8_l16384_id3_1_0_wenable(ram_w8_l16384_id3_1_0_wenable),
    .ram_w8_l16384_id3_1_0_enable(ram_w8_l16384_id3_1_0_enable),
    .ram_w8_l16384_id3_1_1_addr(ram_w8_l16384_id3_1_1_addr),
    .ram_w8_l16384_id3_1_1_rdata(ram_w8_l16384_id3_1_1_rdata),
    .ram_w8_l16384_id3_1_1_wdata(ram_w8_l16384_id3_1_1_wdata),
    .ram_w8_l16384_id3_1_1_wenable(ram_w8_l16384_id3_1_1_wenable),
    .ram_w8_l16384_id3_1_1_enable(ram_w8_l16384_id3_1_1_enable)
  );

  wire [12-1:0] ram_w8_l16384_id3_2_0_addr;
  wire [8-1:0] ram_w8_l16384_id3_2_0_rdata;
  wire [8-1:0] ram_w8_l16384_id3_2_0_wdata;
  wire ram_w8_l16384_id3_2_0_wenable;
  wire ram_w8_l16384_id3_2_0_enable;
  wire [12-1:0] ram_w8_l16384_id3_2_1_addr;
  wire [8-1:0] ram_w8_l16384_id3_2_1_rdata;
  wire [8-1:0] ram_w8_l16384_id3_2_1_wdata;
  wire ram_w8_l16384_id3_2_1_wenable;
  wire ram_w8_l16384_id3_2_1_enable;
  assign ram_w8_l16384_id3_2_0_wdata = 'hx;
  assign ram_w8_l16384_id3_2_0_wenable = 0;

  ram_w8_l16384_id3_2
  inst_ram_w8_l16384_id3_2
  (
    .CLK(CLK),
    .ram_w8_l16384_id3_2_0_addr(ram_w8_l16384_id3_2_0_addr),
    .ram_w8_l16384_id3_2_0_rdata(ram_w8_l16384_id3_2_0_rdata),
    .ram_w8_l16384_id3_2_0_wdata(ram_w8_l16384_id3_2_0_wdata),
    .ram_w8_l16384_id3_2_0_wenable(ram_w8_l16384_id3_2_0_wenable),
    .ram_w8_l16384_id3_2_0_enable(ram_w8_l16384_id3_2_0_enable),
    .ram_w8_l16384_id3_2_1_addr(ram_w8_l16384_id3_2_1_addr),
    .ram_w8_l16384_id3_2_1_rdata(ram_w8_l16384_id3_2_1_rdata),
    .ram_w8_l16384_id3_2_1_wdata(ram_w8_l16384_id3_2_1_wdata),
    .ram_w8_l16384_id3_2_1_wenable(ram_w8_l16384_id3_2_1_wenable),
    .ram_w8_l16384_id3_2_1_enable(ram_w8_l16384_id3_2_1_enable)
  );

  wire [12-1:0] ram_w8_l16384_id3_3_0_addr;
  wire [8-1:0] ram_w8_l16384_id3_3_0_rdata;
  wire [8-1:0] ram_w8_l16384_id3_3_0_wdata;
  wire ram_w8_l16384_id3_3_0_wenable;
  wire ram_w8_l16384_id3_3_0_enable;
  wire [12-1:0] ram_w8_l16384_id3_3_1_addr;
  wire [8-1:0] ram_w8_l16384_id3_3_1_rdata;
  wire [8-1:0] ram_w8_l16384_id3_3_1_wdata;
  wire ram_w8_l16384_id3_3_1_wenable;
  wire ram_w8_l16384_id3_3_1_enable;
  assign ram_w8_l16384_id3_3_0_wdata = 'hx;
  assign ram_w8_l16384_id3_3_0_wenable = 0;

  ram_w8_l16384_id3_3
  inst_ram_w8_l16384_id3_3
  (
    .CLK(CLK),
    .ram_w8_l16384_id3_3_0_addr(ram_w8_l16384_id3_3_0_addr),
    .ram_w8_l16384_id3_3_0_rdata(ram_w8_l16384_id3_3_0_rdata),
    .ram_w8_l16384_id3_3_0_wdata(ram_w8_l16384_id3_3_0_wdata),
    .ram_w8_l16384_id3_3_0_wenable(ram_w8_l16384_id3_3_0_wenable),
    .ram_w8_l16384_id3_3_0_enable(ram_w8_l16384_id3_3_0_enable),
    .ram_w8_l16384_id3_3_1_addr(ram_w8_l16384_id3_3_1_addr),
    .ram_w8_l16384_id3_3_1_rdata(ram_w8_l16384_id3_3_1_rdata),
    .ram_w8_l16384_id3_3_1_wdata(ram_w8_l16384_id3_3_1_wdata),
    .ram_w8_l16384_id3_3_1_wenable(ram_w8_l16384_id3_3_1_wenable),
    .ram_w8_l16384_id3_3_1_enable(ram_w8_l16384_id3_3_1_enable)
  );

  wire [12-1:0] ram_w8_l16384_id4_0_0_addr;
  wire [8-1:0] ram_w8_l16384_id4_0_0_rdata;
  wire [8-1:0] ram_w8_l16384_id4_0_0_wdata;
  wire ram_w8_l16384_id4_0_0_wenable;
  wire ram_w8_l16384_id4_0_0_enable;
  wire [12-1:0] ram_w8_l16384_id4_0_1_addr;
  wire [8-1:0] ram_w8_l16384_id4_0_1_rdata;
  wire [8-1:0] ram_w8_l16384_id4_0_1_wdata;
  wire ram_w8_l16384_id4_0_1_wenable;
  wire ram_w8_l16384_id4_0_1_enable;
  assign ram_w8_l16384_id4_0_0_wdata = 'hx;
  assign ram_w8_l16384_id4_0_0_wenable = 0;

  ram_w8_l16384_id4_0
  inst_ram_w8_l16384_id4_0
  (
    .CLK(CLK),
    .ram_w8_l16384_id4_0_0_addr(ram_w8_l16384_id4_0_0_addr),
    .ram_w8_l16384_id4_0_0_rdata(ram_w8_l16384_id4_0_0_rdata),
    .ram_w8_l16384_id4_0_0_wdata(ram_w8_l16384_id4_0_0_wdata),
    .ram_w8_l16384_id4_0_0_wenable(ram_w8_l16384_id4_0_0_wenable),
    .ram_w8_l16384_id4_0_0_enable(ram_w8_l16384_id4_0_0_enable),
    .ram_w8_l16384_id4_0_1_addr(ram_w8_l16384_id4_0_1_addr),
    .ram_w8_l16384_id4_0_1_rdata(ram_w8_l16384_id4_0_1_rdata),
    .ram_w8_l16384_id4_0_1_wdata(ram_w8_l16384_id4_0_1_wdata),
    .ram_w8_l16384_id4_0_1_wenable(ram_w8_l16384_id4_0_1_wenable),
    .ram_w8_l16384_id4_0_1_enable(ram_w8_l16384_id4_0_1_enable)
  );

  wire [12-1:0] ram_w8_l16384_id4_1_0_addr;
  wire [8-1:0] ram_w8_l16384_id4_1_0_rdata;
  wire [8-1:0] ram_w8_l16384_id4_1_0_wdata;
  wire ram_w8_l16384_id4_1_0_wenable;
  wire ram_w8_l16384_id4_1_0_enable;
  wire [12-1:0] ram_w8_l16384_id4_1_1_addr;
  wire [8-1:0] ram_w8_l16384_id4_1_1_rdata;
  wire [8-1:0] ram_w8_l16384_id4_1_1_wdata;
  wire ram_w8_l16384_id4_1_1_wenable;
  wire ram_w8_l16384_id4_1_1_enable;
  assign ram_w8_l16384_id4_1_0_wdata = 'hx;
  assign ram_w8_l16384_id4_1_0_wenable = 0;

  ram_w8_l16384_id4_1
  inst_ram_w8_l16384_id4_1
  (
    .CLK(CLK),
    .ram_w8_l16384_id4_1_0_addr(ram_w8_l16384_id4_1_0_addr),
    .ram_w8_l16384_id4_1_0_rdata(ram_w8_l16384_id4_1_0_rdata),
    .ram_w8_l16384_id4_1_0_wdata(ram_w8_l16384_id4_1_0_wdata),
    .ram_w8_l16384_id4_1_0_wenable(ram_w8_l16384_id4_1_0_wenable),
    .ram_w8_l16384_id4_1_0_enable(ram_w8_l16384_id4_1_0_enable),
    .ram_w8_l16384_id4_1_1_addr(ram_w8_l16384_id4_1_1_addr),
    .ram_w8_l16384_id4_1_1_rdata(ram_w8_l16384_id4_1_1_rdata),
    .ram_w8_l16384_id4_1_1_wdata(ram_w8_l16384_id4_1_1_wdata),
    .ram_w8_l16384_id4_1_1_wenable(ram_w8_l16384_id4_1_1_wenable),
    .ram_w8_l16384_id4_1_1_enable(ram_w8_l16384_id4_1_1_enable)
  );

  wire [12-1:0] ram_w8_l16384_id4_2_0_addr;
  wire [8-1:0] ram_w8_l16384_id4_2_0_rdata;
  wire [8-1:0] ram_w8_l16384_id4_2_0_wdata;
  wire ram_w8_l16384_id4_2_0_wenable;
  wire ram_w8_l16384_id4_2_0_enable;
  wire [12-1:0] ram_w8_l16384_id4_2_1_addr;
  wire [8-1:0] ram_w8_l16384_id4_2_1_rdata;
  wire [8-1:0] ram_w8_l16384_id4_2_1_wdata;
  wire ram_w8_l16384_id4_2_1_wenable;
  wire ram_w8_l16384_id4_2_1_enable;
  assign ram_w8_l16384_id4_2_0_wdata = 'hx;
  assign ram_w8_l16384_id4_2_0_wenable = 0;

  ram_w8_l16384_id4_2
  inst_ram_w8_l16384_id4_2
  (
    .CLK(CLK),
    .ram_w8_l16384_id4_2_0_addr(ram_w8_l16384_id4_2_0_addr),
    .ram_w8_l16384_id4_2_0_rdata(ram_w8_l16384_id4_2_0_rdata),
    .ram_w8_l16384_id4_2_0_wdata(ram_w8_l16384_id4_2_0_wdata),
    .ram_w8_l16384_id4_2_0_wenable(ram_w8_l16384_id4_2_0_wenable),
    .ram_w8_l16384_id4_2_0_enable(ram_w8_l16384_id4_2_0_enable),
    .ram_w8_l16384_id4_2_1_addr(ram_w8_l16384_id4_2_1_addr),
    .ram_w8_l16384_id4_2_1_rdata(ram_w8_l16384_id4_2_1_rdata),
    .ram_w8_l16384_id4_2_1_wdata(ram_w8_l16384_id4_2_1_wdata),
    .ram_w8_l16384_id4_2_1_wenable(ram_w8_l16384_id4_2_1_wenable),
    .ram_w8_l16384_id4_2_1_enable(ram_w8_l16384_id4_2_1_enable)
  );

  wire [12-1:0] ram_w8_l16384_id4_3_0_addr;
  wire [8-1:0] ram_w8_l16384_id4_3_0_rdata;
  wire [8-1:0] ram_w8_l16384_id4_3_0_wdata;
  wire ram_w8_l16384_id4_3_0_wenable;
  wire ram_w8_l16384_id4_3_0_enable;
  wire [12-1:0] ram_w8_l16384_id4_3_1_addr;
  wire [8-1:0] ram_w8_l16384_id4_3_1_rdata;
  wire [8-1:0] ram_w8_l16384_id4_3_1_wdata;
  wire ram_w8_l16384_id4_3_1_wenable;
  wire ram_w8_l16384_id4_3_1_enable;
  assign ram_w8_l16384_id4_3_0_wdata = 'hx;
  assign ram_w8_l16384_id4_3_0_wenable = 0;

  ram_w8_l16384_id4_3
  inst_ram_w8_l16384_id4_3
  (
    .CLK(CLK),
    .ram_w8_l16384_id4_3_0_addr(ram_w8_l16384_id4_3_0_addr),
    .ram_w8_l16384_id4_3_0_rdata(ram_w8_l16384_id4_3_0_rdata),
    .ram_w8_l16384_id4_3_0_wdata(ram_w8_l16384_id4_3_0_wdata),
    .ram_w8_l16384_id4_3_0_wenable(ram_w8_l16384_id4_3_0_wenable),
    .ram_w8_l16384_id4_3_0_enable(ram_w8_l16384_id4_3_0_enable),
    .ram_w8_l16384_id4_3_1_addr(ram_w8_l16384_id4_3_1_addr),
    .ram_w8_l16384_id4_3_1_rdata(ram_w8_l16384_id4_3_1_rdata),
    .ram_w8_l16384_id4_3_1_wdata(ram_w8_l16384_id4_3_1_wdata),
    .ram_w8_l16384_id4_3_1_wenable(ram_w8_l16384_id4_3_1_wenable),
    .ram_w8_l16384_id4_3_1_enable(ram_w8_l16384_id4_3_1_enable)
  );

  wire [12-1:0] ram_w8_l16384_id5_0_0_addr;
  wire [8-1:0] ram_w8_l16384_id5_0_0_rdata;
  wire [8-1:0] ram_w8_l16384_id5_0_0_wdata;
  wire ram_w8_l16384_id5_0_0_wenable;
  wire ram_w8_l16384_id5_0_0_enable;
  wire [12-1:0] ram_w8_l16384_id5_0_1_addr;
  wire [8-1:0] ram_w8_l16384_id5_0_1_rdata;
  wire [8-1:0] ram_w8_l16384_id5_0_1_wdata;
  wire ram_w8_l16384_id5_0_1_wenable;
  wire ram_w8_l16384_id5_0_1_enable;
  assign ram_w8_l16384_id5_0_0_wdata = 'hx;
  assign ram_w8_l16384_id5_0_0_wenable = 0;

  ram_w8_l16384_id5_0
  inst_ram_w8_l16384_id5_0
  (
    .CLK(CLK),
    .ram_w8_l16384_id5_0_0_addr(ram_w8_l16384_id5_0_0_addr),
    .ram_w8_l16384_id5_0_0_rdata(ram_w8_l16384_id5_0_0_rdata),
    .ram_w8_l16384_id5_0_0_wdata(ram_w8_l16384_id5_0_0_wdata),
    .ram_w8_l16384_id5_0_0_wenable(ram_w8_l16384_id5_0_0_wenable),
    .ram_w8_l16384_id5_0_0_enable(ram_w8_l16384_id5_0_0_enable),
    .ram_w8_l16384_id5_0_1_addr(ram_w8_l16384_id5_0_1_addr),
    .ram_w8_l16384_id5_0_1_rdata(ram_w8_l16384_id5_0_1_rdata),
    .ram_w8_l16384_id5_0_1_wdata(ram_w8_l16384_id5_0_1_wdata),
    .ram_w8_l16384_id5_0_1_wenable(ram_w8_l16384_id5_0_1_wenable),
    .ram_w8_l16384_id5_0_1_enable(ram_w8_l16384_id5_0_1_enable)
  );

  wire [12-1:0] ram_w8_l16384_id5_1_0_addr;
  wire [8-1:0] ram_w8_l16384_id5_1_0_rdata;
  wire [8-1:0] ram_w8_l16384_id5_1_0_wdata;
  wire ram_w8_l16384_id5_1_0_wenable;
  wire ram_w8_l16384_id5_1_0_enable;
  wire [12-1:0] ram_w8_l16384_id5_1_1_addr;
  wire [8-1:0] ram_w8_l16384_id5_1_1_rdata;
  wire [8-1:0] ram_w8_l16384_id5_1_1_wdata;
  wire ram_w8_l16384_id5_1_1_wenable;
  wire ram_w8_l16384_id5_1_1_enable;
  assign ram_w8_l16384_id5_1_0_wdata = 'hx;
  assign ram_w8_l16384_id5_1_0_wenable = 0;

  ram_w8_l16384_id5_1
  inst_ram_w8_l16384_id5_1
  (
    .CLK(CLK),
    .ram_w8_l16384_id5_1_0_addr(ram_w8_l16384_id5_1_0_addr),
    .ram_w8_l16384_id5_1_0_rdata(ram_w8_l16384_id5_1_0_rdata),
    .ram_w8_l16384_id5_1_0_wdata(ram_w8_l16384_id5_1_0_wdata),
    .ram_w8_l16384_id5_1_0_wenable(ram_w8_l16384_id5_1_0_wenable),
    .ram_w8_l16384_id5_1_0_enable(ram_w8_l16384_id5_1_0_enable),
    .ram_w8_l16384_id5_1_1_addr(ram_w8_l16384_id5_1_1_addr),
    .ram_w8_l16384_id5_1_1_rdata(ram_w8_l16384_id5_1_1_rdata),
    .ram_w8_l16384_id5_1_1_wdata(ram_w8_l16384_id5_1_1_wdata),
    .ram_w8_l16384_id5_1_1_wenable(ram_w8_l16384_id5_1_1_wenable),
    .ram_w8_l16384_id5_1_1_enable(ram_w8_l16384_id5_1_1_enable)
  );

  wire [12-1:0] ram_w8_l16384_id5_2_0_addr;
  wire [8-1:0] ram_w8_l16384_id5_2_0_rdata;
  wire [8-1:0] ram_w8_l16384_id5_2_0_wdata;
  wire ram_w8_l16384_id5_2_0_wenable;
  wire ram_w8_l16384_id5_2_0_enable;
  wire [12-1:0] ram_w8_l16384_id5_2_1_addr;
  wire [8-1:0] ram_w8_l16384_id5_2_1_rdata;
  wire [8-1:0] ram_w8_l16384_id5_2_1_wdata;
  wire ram_w8_l16384_id5_2_1_wenable;
  wire ram_w8_l16384_id5_2_1_enable;
  assign ram_w8_l16384_id5_2_0_wdata = 'hx;
  assign ram_w8_l16384_id5_2_0_wenable = 0;

  ram_w8_l16384_id5_2
  inst_ram_w8_l16384_id5_2
  (
    .CLK(CLK),
    .ram_w8_l16384_id5_2_0_addr(ram_w8_l16384_id5_2_0_addr),
    .ram_w8_l16384_id5_2_0_rdata(ram_w8_l16384_id5_2_0_rdata),
    .ram_w8_l16384_id5_2_0_wdata(ram_w8_l16384_id5_2_0_wdata),
    .ram_w8_l16384_id5_2_0_wenable(ram_w8_l16384_id5_2_0_wenable),
    .ram_w8_l16384_id5_2_0_enable(ram_w8_l16384_id5_2_0_enable),
    .ram_w8_l16384_id5_2_1_addr(ram_w8_l16384_id5_2_1_addr),
    .ram_w8_l16384_id5_2_1_rdata(ram_w8_l16384_id5_2_1_rdata),
    .ram_w8_l16384_id5_2_1_wdata(ram_w8_l16384_id5_2_1_wdata),
    .ram_w8_l16384_id5_2_1_wenable(ram_w8_l16384_id5_2_1_wenable),
    .ram_w8_l16384_id5_2_1_enable(ram_w8_l16384_id5_2_1_enable)
  );

  wire [12-1:0] ram_w8_l16384_id5_3_0_addr;
  wire [8-1:0] ram_w8_l16384_id5_3_0_rdata;
  wire [8-1:0] ram_w8_l16384_id5_3_0_wdata;
  wire ram_w8_l16384_id5_3_0_wenable;
  wire ram_w8_l16384_id5_3_0_enable;
  wire [12-1:0] ram_w8_l16384_id5_3_1_addr;
  wire [8-1:0] ram_w8_l16384_id5_3_1_rdata;
  wire [8-1:0] ram_w8_l16384_id5_3_1_wdata;
  wire ram_w8_l16384_id5_3_1_wenable;
  wire ram_w8_l16384_id5_3_1_enable;
  assign ram_w8_l16384_id5_3_0_wdata = 'hx;
  assign ram_w8_l16384_id5_3_0_wenable = 0;

  ram_w8_l16384_id5_3
  inst_ram_w8_l16384_id5_3
  (
    .CLK(CLK),
    .ram_w8_l16384_id5_3_0_addr(ram_w8_l16384_id5_3_0_addr),
    .ram_w8_l16384_id5_3_0_rdata(ram_w8_l16384_id5_3_0_rdata),
    .ram_w8_l16384_id5_3_0_wdata(ram_w8_l16384_id5_3_0_wdata),
    .ram_w8_l16384_id5_3_0_wenable(ram_w8_l16384_id5_3_0_wenable),
    .ram_w8_l16384_id5_3_0_enable(ram_w8_l16384_id5_3_0_enable),
    .ram_w8_l16384_id5_3_1_addr(ram_w8_l16384_id5_3_1_addr),
    .ram_w8_l16384_id5_3_1_rdata(ram_w8_l16384_id5_3_1_rdata),
    .ram_w8_l16384_id5_3_1_wdata(ram_w8_l16384_id5_3_1_wdata),
    .ram_w8_l16384_id5_3_1_wenable(ram_w8_l16384_id5_3_1_wenable),
    .ram_w8_l16384_id5_3_1_enable(ram_w8_l16384_id5_3_1_enable)
  );

  wire [12-1:0] ram_w8_l16384_id6_0_0_addr;
  wire [8-1:0] ram_w8_l16384_id6_0_0_rdata;
  wire [8-1:0] ram_w8_l16384_id6_0_0_wdata;
  wire ram_w8_l16384_id6_0_0_wenable;
  wire ram_w8_l16384_id6_0_0_enable;
  wire [12-1:0] ram_w8_l16384_id6_0_1_addr;
  wire [8-1:0] ram_w8_l16384_id6_0_1_rdata;
  wire [8-1:0] ram_w8_l16384_id6_0_1_wdata;
  wire ram_w8_l16384_id6_0_1_wenable;
  wire ram_w8_l16384_id6_0_1_enable;
  assign ram_w8_l16384_id6_0_0_wdata = 'hx;
  assign ram_w8_l16384_id6_0_0_wenable = 0;

  ram_w8_l16384_id6_0
  inst_ram_w8_l16384_id6_0
  (
    .CLK(CLK),
    .ram_w8_l16384_id6_0_0_addr(ram_w8_l16384_id6_0_0_addr),
    .ram_w8_l16384_id6_0_0_rdata(ram_w8_l16384_id6_0_0_rdata),
    .ram_w8_l16384_id6_0_0_wdata(ram_w8_l16384_id6_0_0_wdata),
    .ram_w8_l16384_id6_0_0_wenable(ram_w8_l16384_id6_0_0_wenable),
    .ram_w8_l16384_id6_0_0_enable(ram_w8_l16384_id6_0_0_enable),
    .ram_w8_l16384_id6_0_1_addr(ram_w8_l16384_id6_0_1_addr),
    .ram_w8_l16384_id6_0_1_rdata(ram_w8_l16384_id6_0_1_rdata),
    .ram_w8_l16384_id6_0_1_wdata(ram_w8_l16384_id6_0_1_wdata),
    .ram_w8_l16384_id6_0_1_wenable(ram_w8_l16384_id6_0_1_wenable),
    .ram_w8_l16384_id6_0_1_enable(ram_w8_l16384_id6_0_1_enable)
  );

  wire [12-1:0] ram_w8_l16384_id6_1_0_addr;
  wire [8-1:0] ram_w8_l16384_id6_1_0_rdata;
  wire [8-1:0] ram_w8_l16384_id6_1_0_wdata;
  wire ram_w8_l16384_id6_1_0_wenable;
  wire ram_w8_l16384_id6_1_0_enable;
  wire [12-1:0] ram_w8_l16384_id6_1_1_addr;
  wire [8-1:0] ram_w8_l16384_id6_1_1_rdata;
  wire [8-1:0] ram_w8_l16384_id6_1_1_wdata;
  wire ram_w8_l16384_id6_1_1_wenable;
  wire ram_w8_l16384_id6_1_1_enable;
  assign ram_w8_l16384_id6_1_0_wdata = 'hx;
  assign ram_w8_l16384_id6_1_0_wenable = 0;

  ram_w8_l16384_id6_1
  inst_ram_w8_l16384_id6_1
  (
    .CLK(CLK),
    .ram_w8_l16384_id6_1_0_addr(ram_w8_l16384_id6_1_0_addr),
    .ram_w8_l16384_id6_1_0_rdata(ram_w8_l16384_id6_1_0_rdata),
    .ram_w8_l16384_id6_1_0_wdata(ram_w8_l16384_id6_1_0_wdata),
    .ram_w8_l16384_id6_1_0_wenable(ram_w8_l16384_id6_1_0_wenable),
    .ram_w8_l16384_id6_1_0_enable(ram_w8_l16384_id6_1_0_enable),
    .ram_w8_l16384_id6_1_1_addr(ram_w8_l16384_id6_1_1_addr),
    .ram_w8_l16384_id6_1_1_rdata(ram_w8_l16384_id6_1_1_rdata),
    .ram_w8_l16384_id6_1_1_wdata(ram_w8_l16384_id6_1_1_wdata),
    .ram_w8_l16384_id6_1_1_wenable(ram_w8_l16384_id6_1_1_wenable),
    .ram_w8_l16384_id6_1_1_enable(ram_w8_l16384_id6_1_1_enable)
  );

  wire [12-1:0] ram_w8_l16384_id6_2_0_addr;
  wire [8-1:0] ram_w8_l16384_id6_2_0_rdata;
  wire [8-1:0] ram_w8_l16384_id6_2_0_wdata;
  wire ram_w8_l16384_id6_2_0_wenable;
  wire ram_w8_l16384_id6_2_0_enable;
  wire [12-1:0] ram_w8_l16384_id6_2_1_addr;
  wire [8-1:0] ram_w8_l16384_id6_2_1_rdata;
  wire [8-1:0] ram_w8_l16384_id6_2_1_wdata;
  wire ram_w8_l16384_id6_2_1_wenable;
  wire ram_w8_l16384_id6_2_1_enable;
  assign ram_w8_l16384_id6_2_0_wdata = 'hx;
  assign ram_w8_l16384_id6_2_0_wenable = 0;

  ram_w8_l16384_id6_2
  inst_ram_w8_l16384_id6_2
  (
    .CLK(CLK),
    .ram_w8_l16384_id6_2_0_addr(ram_w8_l16384_id6_2_0_addr),
    .ram_w8_l16384_id6_2_0_rdata(ram_w8_l16384_id6_2_0_rdata),
    .ram_w8_l16384_id6_2_0_wdata(ram_w8_l16384_id6_2_0_wdata),
    .ram_w8_l16384_id6_2_0_wenable(ram_w8_l16384_id6_2_0_wenable),
    .ram_w8_l16384_id6_2_0_enable(ram_w8_l16384_id6_2_0_enable),
    .ram_w8_l16384_id6_2_1_addr(ram_w8_l16384_id6_2_1_addr),
    .ram_w8_l16384_id6_2_1_rdata(ram_w8_l16384_id6_2_1_rdata),
    .ram_w8_l16384_id6_2_1_wdata(ram_w8_l16384_id6_2_1_wdata),
    .ram_w8_l16384_id6_2_1_wenable(ram_w8_l16384_id6_2_1_wenable),
    .ram_w8_l16384_id6_2_1_enable(ram_w8_l16384_id6_2_1_enable)
  );

  wire [12-1:0] ram_w8_l16384_id6_3_0_addr;
  wire [8-1:0] ram_w8_l16384_id6_3_0_rdata;
  wire [8-1:0] ram_w8_l16384_id6_3_0_wdata;
  wire ram_w8_l16384_id6_3_0_wenable;
  wire ram_w8_l16384_id6_3_0_enable;
  wire [12-1:0] ram_w8_l16384_id6_3_1_addr;
  wire [8-1:0] ram_w8_l16384_id6_3_1_rdata;
  wire [8-1:0] ram_w8_l16384_id6_3_1_wdata;
  wire ram_w8_l16384_id6_3_1_wenable;
  wire ram_w8_l16384_id6_3_1_enable;
  assign ram_w8_l16384_id6_3_0_wdata = 'hx;
  assign ram_w8_l16384_id6_3_0_wenable = 0;

  ram_w8_l16384_id6_3
  inst_ram_w8_l16384_id6_3
  (
    .CLK(CLK),
    .ram_w8_l16384_id6_3_0_addr(ram_w8_l16384_id6_3_0_addr),
    .ram_w8_l16384_id6_3_0_rdata(ram_w8_l16384_id6_3_0_rdata),
    .ram_w8_l16384_id6_3_0_wdata(ram_w8_l16384_id6_3_0_wdata),
    .ram_w8_l16384_id6_3_0_wenable(ram_w8_l16384_id6_3_0_wenable),
    .ram_w8_l16384_id6_3_0_enable(ram_w8_l16384_id6_3_0_enable),
    .ram_w8_l16384_id6_3_1_addr(ram_w8_l16384_id6_3_1_addr),
    .ram_w8_l16384_id6_3_1_rdata(ram_w8_l16384_id6_3_1_rdata),
    .ram_w8_l16384_id6_3_1_wdata(ram_w8_l16384_id6_3_1_wdata),
    .ram_w8_l16384_id6_3_1_wenable(ram_w8_l16384_id6_3_1_wenable),
    .ram_w8_l16384_id6_3_1_enable(ram_w8_l16384_id6_3_1_enable)
  );

  wire [12-1:0] ram_w8_l16384_id7_0_0_addr;
  wire [8-1:0] ram_w8_l16384_id7_0_0_rdata;
  wire [8-1:0] ram_w8_l16384_id7_0_0_wdata;
  wire ram_w8_l16384_id7_0_0_wenable;
  wire ram_w8_l16384_id7_0_0_enable;
  wire [12-1:0] ram_w8_l16384_id7_0_1_addr;
  wire [8-1:0] ram_w8_l16384_id7_0_1_rdata;
  wire [8-1:0] ram_w8_l16384_id7_0_1_wdata;
  wire ram_w8_l16384_id7_0_1_wenable;
  wire ram_w8_l16384_id7_0_1_enable;
  assign ram_w8_l16384_id7_0_0_wdata = 'hx;
  assign ram_w8_l16384_id7_0_0_wenable = 0;

  ram_w8_l16384_id7_0
  inst_ram_w8_l16384_id7_0
  (
    .CLK(CLK),
    .ram_w8_l16384_id7_0_0_addr(ram_w8_l16384_id7_0_0_addr),
    .ram_w8_l16384_id7_0_0_rdata(ram_w8_l16384_id7_0_0_rdata),
    .ram_w8_l16384_id7_0_0_wdata(ram_w8_l16384_id7_0_0_wdata),
    .ram_w8_l16384_id7_0_0_wenable(ram_w8_l16384_id7_0_0_wenable),
    .ram_w8_l16384_id7_0_0_enable(ram_w8_l16384_id7_0_0_enable),
    .ram_w8_l16384_id7_0_1_addr(ram_w8_l16384_id7_0_1_addr),
    .ram_w8_l16384_id7_0_1_rdata(ram_w8_l16384_id7_0_1_rdata),
    .ram_w8_l16384_id7_0_1_wdata(ram_w8_l16384_id7_0_1_wdata),
    .ram_w8_l16384_id7_0_1_wenable(ram_w8_l16384_id7_0_1_wenable),
    .ram_w8_l16384_id7_0_1_enable(ram_w8_l16384_id7_0_1_enable)
  );

  wire [12-1:0] ram_w8_l16384_id7_1_0_addr;
  wire [8-1:0] ram_w8_l16384_id7_1_0_rdata;
  wire [8-1:0] ram_w8_l16384_id7_1_0_wdata;
  wire ram_w8_l16384_id7_1_0_wenable;
  wire ram_w8_l16384_id7_1_0_enable;
  wire [12-1:0] ram_w8_l16384_id7_1_1_addr;
  wire [8-1:0] ram_w8_l16384_id7_1_1_rdata;
  wire [8-1:0] ram_w8_l16384_id7_1_1_wdata;
  wire ram_w8_l16384_id7_1_1_wenable;
  wire ram_w8_l16384_id7_1_1_enable;
  assign ram_w8_l16384_id7_1_0_wdata = 'hx;
  assign ram_w8_l16384_id7_1_0_wenable = 0;

  ram_w8_l16384_id7_1
  inst_ram_w8_l16384_id7_1
  (
    .CLK(CLK),
    .ram_w8_l16384_id7_1_0_addr(ram_w8_l16384_id7_1_0_addr),
    .ram_w8_l16384_id7_1_0_rdata(ram_w8_l16384_id7_1_0_rdata),
    .ram_w8_l16384_id7_1_0_wdata(ram_w8_l16384_id7_1_0_wdata),
    .ram_w8_l16384_id7_1_0_wenable(ram_w8_l16384_id7_1_0_wenable),
    .ram_w8_l16384_id7_1_0_enable(ram_w8_l16384_id7_1_0_enable),
    .ram_w8_l16384_id7_1_1_addr(ram_w8_l16384_id7_1_1_addr),
    .ram_w8_l16384_id7_1_1_rdata(ram_w8_l16384_id7_1_1_rdata),
    .ram_w8_l16384_id7_1_1_wdata(ram_w8_l16384_id7_1_1_wdata),
    .ram_w8_l16384_id7_1_1_wenable(ram_w8_l16384_id7_1_1_wenable),
    .ram_w8_l16384_id7_1_1_enable(ram_w8_l16384_id7_1_1_enable)
  );

  wire [12-1:0] ram_w8_l16384_id7_2_0_addr;
  wire [8-1:0] ram_w8_l16384_id7_2_0_rdata;
  wire [8-1:0] ram_w8_l16384_id7_2_0_wdata;
  wire ram_w8_l16384_id7_2_0_wenable;
  wire ram_w8_l16384_id7_2_0_enable;
  wire [12-1:0] ram_w8_l16384_id7_2_1_addr;
  wire [8-1:0] ram_w8_l16384_id7_2_1_rdata;
  wire [8-1:0] ram_w8_l16384_id7_2_1_wdata;
  wire ram_w8_l16384_id7_2_1_wenable;
  wire ram_w8_l16384_id7_2_1_enable;
  assign ram_w8_l16384_id7_2_0_wdata = 'hx;
  assign ram_w8_l16384_id7_2_0_wenable = 0;

  ram_w8_l16384_id7_2
  inst_ram_w8_l16384_id7_2
  (
    .CLK(CLK),
    .ram_w8_l16384_id7_2_0_addr(ram_w8_l16384_id7_2_0_addr),
    .ram_w8_l16384_id7_2_0_rdata(ram_w8_l16384_id7_2_0_rdata),
    .ram_w8_l16384_id7_2_0_wdata(ram_w8_l16384_id7_2_0_wdata),
    .ram_w8_l16384_id7_2_0_wenable(ram_w8_l16384_id7_2_0_wenable),
    .ram_w8_l16384_id7_2_0_enable(ram_w8_l16384_id7_2_0_enable),
    .ram_w8_l16384_id7_2_1_addr(ram_w8_l16384_id7_2_1_addr),
    .ram_w8_l16384_id7_2_1_rdata(ram_w8_l16384_id7_2_1_rdata),
    .ram_w8_l16384_id7_2_1_wdata(ram_w8_l16384_id7_2_1_wdata),
    .ram_w8_l16384_id7_2_1_wenable(ram_w8_l16384_id7_2_1_wenable),
    .ram_w8_l16384_id7_2_1_enable(ram_w8_l16384_id7_2_1_enable)
  );

  wire [12-1:0] ram_w8_l16384_id7_3_0_addr;
  wire [8-1:0] ram_w8_l16384_id7_3_0_rdata;
  wire [8-1:0] ram_w8_l16384_id7_3_0_wdata;
  wire ram_w8_l16384_id7_3_0_wenable;
  wire ram_w8_l16384_id7_3_0_enable;
  wire [12-1:0] ram_w8_l16384_id7_3_1_addr;
  wire [8-1:0] ram_w8_l16384_id7_3_1_rdata;
  wire [8-1:0] ram_w8_l16384_id7_3_1_wdata;
  wire ram_w8_l16384_id7_3_1_wenable;
  wire ram_w8_l16384_id7_3_1_enable;
  assign ram_w8_l16384_id7_3_0_wdata = 'hx;
  assign ram_w8_l16384_id7_3_0_wenable = 0;

  ram_w8_l16384_id7_3
  inst_ram_w8_l16384_id7_3
  (
    .CLK(CLK),
    .ram_w8_l16384_id7_3_0_addr(ram_w8_l16384_id7_3_0_addr),
    .ram_w8_l16384_id7_3_0_rdata(ram_w8_l16384_id7_3_0_rdata),
    .ram_w8_l16384_id7_3_0_wdata(ram_w8_l16384_id7_3_0_wdata),
    .ram_w8_l16384_id7_3_0_wenable(ram_w8_l16384_id7_3_0_wenable),
    .ram_w8_l16384_id7_3_0_enable(ram_w8_l16384_id7_3_0_enable),
    .ram_w8_l16384_id7_3_1_addr(ram_w8_l16384_id7_3_1_addr),
    .ram_w8_l16384_id7_3_1_rdata(ram_w8_l16384_id7_3_1_rdata),
    .ram_w8_l16384_id7_3_1_wdata(ram_w8_l16384_id7_3_1_wdata),
    .ram_w8_l16384_id7_3_1_wenable(ram_w8_l16384_id7_3_1_wenable),
    .ram_w8_l16384_id7_3_1_enable(ram_w8_l16384_id7_3_1_enable)
  );

  wire [12-1:0] ram_w8_l16384_id8_0_0_addr;
  wire [8-1:0] ram_w8_l16384_id8_0_0_rdata;
  wire [8-1:0] ram_w8_l16384_id8_0_0_wdata;
  wire ram_w8_l16384_id8_0_0_wenable;
  wire ram_w8_l16384_id8_0_0_enable;
  wire [12-1:0] ram_w8_l16384_id8_0_1_addr;
  wire [8-1:0] ram_w8_l16384_id8_0_1_rdata;
  wire [8-1:0] ram_w8_l16384_id8_0_1_wdata;
  wire ram_w8_l16384_id8_0_1_wenable;
  wire ram_w8_l16384_id8_0_1_enable;
  assign ram_w8_l16384_id8_0_0_wdata = 'hx;
  assign ram_w8_l16384_id8_0_0_wenable = 0;

  ram_w8_l16384_id8_0
  inst_ram_w8_l16384_id8_0
  (
    .CLK(CLK),
    .ram_w8_l16384_id8_0_0_addr(ram_w8_l16384_id8_0_0_addr),
    .ram_w8_l16384_id8_0_0_rdata(ram_w8_l16384_id8_0_0_rdata),
    .ram_w8_l16384_id8_0_0_wdata(ram_w8_l16384_id8_0_0_wdata),
    .ram_w8_l16384_id8_0_0_wenable(ram_w8_l16384_id8_0_0_wenable),
    .ram_w8_l16384_id8_0_0_enable(ram_w8_l16384_id8_0_0_enable),
    .ram_w8_l16384_id8_0_1_addr(ram_w8_l16384_id8_0_1_addr),
    .ram_w8_l16384_id8_0_1_rdata(ram_w8_l16384_id8_0_1_rdata),
    .ram_w8_l16384_id8_0_1_wdata(ram_w8_l16384_id8_0_1_wdata),
    .ram_w8_l16384_id8_0_1_wenable(ram_w8_l16384_id8_0_1_wenable),
    .ram_w8_l16384_id8_0_1_enable(ram_w8_l16384_id8_0_1_enable)
  );

  wire [12-1:0] ram_w8_l16384_id8_1_0_addr;
  wire [8-1:0] ram_w8_l16384_id8_1_0_rdata;
  wire [8-1:0] ram_w8_l16384_id8_1_0_wdata;
  wire ram_w8_l16384_id8_1_0_wenable;
  wire ram_w8_l16384_id8_1_0_enable;
  wire [12-1:0] ram_w8_l16384_id8_1_1_addr;
  wire [8-1:0] ram_w8_l16384_id8_1_1_rdata;
  wire [8-1:0] ram_w8_l16384_id8_1_1_wdata;
  wire ram_w8_l16384_id8_1_1_wenable;
  wire ram_w8_l16384_id8_1_1_enable;
  assign ram_w8_l16384_id8_1_0_wdata = 'hx;
  assign ram_w8_l16384_id8_1_0_wenable = 0;

  ram_w8_l16384_id8_1
  inst_ram_w8_l16384_id8_1
  (
    .CLK(CLK),
    .ram_w8_l16384_id8_1_0_addr(ram_w8_l16384_id8_1_0_addr),
    .ram_w8_l16384_id8_1_0_rdata(ram_w8_l16384_id8_1_0_rdata),
    .ram_w8_l16384_id8_1_0_wdata(ram_w8_l16384_id8_1_0_wdata),
    .ram_w8_l16384_id8_1_0_wenable(ram_w8_l16384_id8_1_0_wenable),
    .ram_w8_l16384_id8_1_0_enable(ram_w8_l16384_id8_1_0_enable),
    .ram_w8_l16384_id8_1_1_addr(ram_w8_l16384_id8_1_1_addr),
    .ram_w8_l16384_id8_1_1_rdata(ram_w8_l16384_id8_1_1_rdata),
    .ram_w8_l16384_id8_1_1_wdata(ram_w8_l16384_id8_1_1_wdata),
    .ram_w8_l16384_id8_1_1_wenable(ram_w8_l16384_id8_1_1_wenable),
    .ram_w8_l16384_id8_1_1_enable(ram_w8_l16384_id8_1_1_enable)
  );

  wire [12-1:0] ram_w8_l16384_id8_2_0_addr;
  wire [8-1:0] ram_w8_l16384_id8_2_0_rdata;
  wire [8-1:0] ram_w8_l16384_id8_2_0_wdata;
  wire ram_w8_l16384_id8_2_0_wenable;
  wire ram_w8_l16384_id8_2_0_enable;
  wire [12-1:0] ram_w8_l16384_id8_2_1_addr;
  wire [8-1:0] ram_w8_l16384_id8_2_1_rdata;
  wire [8-1:0] ram_w8_l16384_id8_2_1_wdata;
  wire ram_w8_l16384_id8_2_1_wenable;
  wire ram_w8_l16384_id8_2_1_enable;
  assign ram_w8_l16384_id8_2_0_wdata = 'hx;
  assign ram_w8_l16384_id8_2_0_wenable = 0;

  ram_w8_l16384_id8_2
  inst_ram_w8_l16384_id8_2
  (
    .CLK(CLK),
    .ram_w8_l16384_id8_2_0_addr(ram_w8_l16384_id8_2_0_addr),
    .ram_w8_l16384_id8_2_0_rdata(ram_w8_l16384_id8_2_0_rdata),
    .ram_w8_l16384_id8_2_0_wdata(ram_w8_l16384_id8_2_0_wdata),
    .ram_w8_l16384_id8_2_0_wenable(ram_w8_l16384_id8_2_0_wenable),
    .ram_w8_l16384_id8_2_0_enable(ram_w8_l16384_id8_2_0_enable),
    .ram_w8_l16384_id8_2_1_addr(ram_w8_l16384_id8_2_1_addr),
    .ram_w8_l16384_id8_2_1_rdata(ram_w8_l16384_id8_2_1_rdata),
    .ram_w8_l16384_id8_2_1_wdata(ram_w8_l16384_id8_2_1_wdata),
    .ram_w8_l16384_id8_2_1_wenable(ram_w8_l16384_id8_2_1_wenable),
    .ram_w8_l16384_id8_2_1_enable(ram_w8_l16384_id8_2_1_enable)
  );

  wire [12-1:0] ram_w8_l16384_id8_3_0_addr;
  wire [8-1:0] ram_w8_l16384_id8_3_0_rdata;
  wire [8-1:0] ram_w8_l16384_id8_3_0_wdata;
  wire ram_w8_l16384_id8_3_0_wenable;
  wire ram_w8_l16384_id8_3_0_enable;
  wire [12-1:0] ram_w8_l16384_id8_3_1_addr;
  wire [8-1:0] ram_w8_l16384_id8_3_1_rdata;
  wire [8-1:0] ram_w8_l16384_id8_3_1_wdata;
  wire ram_w8_l16384_id8_3_1_wenable;
  wire ram_w8_l16384_id8_3_1_enable;
  assign ram_w8_l16384_id8_3_0_wdata = 'hx;
  assign ram_w8_l16384_id8_3_0_wenable = 0;

  ram_w8_l16384_id8_3
  inst_ram_w8_l16384_id8_3
  (
    .CLK(CLK),
    .ram_w8_l16384_id8_3_0_addr(ram_w8_l16384_id8_3_0_addr),
    .ram_w8_l16384_id8_3_0_rdata(ram_w8_l16384_id8_3_0_rdata),
    .ram_w8_l16384_id8_3_0_wdata(ram_w8_l16384_id8_3_0_wdata),
    .ram_w8_l16384_id8_3_0_wenable(ram_w8_l16384_id8_3_0_wenable),
    .ram_w8_l16384_id8_3_0_enable(ram_w8_l16384_id8_3_0_enable),
    .ram_w8_l16384_id8_3_1_addr(ram_w8_l16384_id8_3_1_addr),
    .ram_w8_l16384_id8_3_1_rdata(ram_w8_l16384_id8_3_1_rdata),
    .ram_w8_l16384_id8_3_1_wdata(ram_w8_l16384_id8_3_1_wdata),
    .ram_w8_l16384_id8_3_1_wenable(ram_w8_l16384_id8_3_1_wenable),
    .ram_w8_l16384_id8_3_1_enable(ram_w8_l16384_id8_3_1_enable)
  );

  wire [12-1:0] ram_w32_l4096_id0_0_addr;
  wire [32-1:0] ram_w32_l4096_id0_0_rdata;
  wire [32-1:0] ram_w32_l4096_id0_0_wdata;
  wire ram_w32_l4096_id0_0_wenable;
  wire ram_w32_l4096_id0_0_enable;
  wire [12-1:0] ram_w32_l4096_id0_1_addr;
  wire [32-1:0] ram_w32_l4096_id0_1_rdata;
  wire [32-1:0] ram_w32_l4096_id0_1_wdata;
  wire ram_w32_l4096_id0_1_wenable;
  wire ram_w32_l4096_id0_1_enable;
  assign ram_w32_l4096_id0_0_wdata = 'hx;
  assign ram_w32_l4096_id0_0_wenable = 0;

  ram_w32_l4096_id0
  inst_ram_w32_l4096_id0
  (
    .CLK(CLK),
    .ram_w32_l4096_id0_0_addr(ram_w32_l4096_id0_0_addr),
    .ram_w32_l4096_id0_0_rdata(ram_w32_l4096_id0_0_rdata),
    .ram_w32_l4096_id0_0_wdata(ram_w32_l4096_id0_0_wdata),
    .ram_w32_l4096_id0_0_wenable(ram_w32_l4096_id0_0_wenable),
    .ram_w32_l4096_id0_0_enable(ram_w32_l4096_id0_0_enable),
    .ram_w32_l4096_id0_1_addr(ram_w32_l4096_id0_1_addr),
    .ram_w32_l4096_id0_1_rdata(ram_w32_l4096_id0_1_rdata),
    .ram_w32_l4096_id0_1_wdata(ram_w32_l4096_id0_1_wdata),
    .ram_w32_l4096_id0_1_wenable(ram_w32_l4096_id0_1_wenable),
    .ram_w32_l4096_id0_1_enable(ram_w32_l4096_id0_1_enable)
  );

  wire [10-1:0] ram_w8_l4096_id0_0_0_addr;
  wire [8-1:0] ram_w8_l4096_id0_0_0_rdata;
  wire [8-1:0] ram_w8_l4096_id0_0_0_wdata;
  wire ram_w8_l4096_id0_0_0_wenable;
  wire ram_w8_l4096_id0_0_0_enable;
  wire [10-1:0] ram_w8_l4096_id0_0_1_addr;
  wire [8-1:0] ram_w8_l4096_id0_0_1_rdata;
  wire [8-1:0] ram_w8_l4096_id0_0_1_wdata;
  wire ram_w8_l4096_id0_0_1_wenable;
  wire ram_w8_l4096_id0_0_1_enable;
  assign ram_w8_l4096_id0_0_0_wdata = 'hx;
  assign ram_w8_l4096_id0_0_0_wenable = 0;

  ram_w8_l4096_id0_0
  inst_ram_w8_l4096_id0_0
  (
    .CLK(CLK),
    .ram_w8_l4096_id0_0_0_addr(ram_w8_l4096_id0_0_0_addr),
    .ram_w8_l4096_id0_0_0_rdata(ram_w8_l4096_id0_0_0_rdata),
    .ram_w8_l4096_id0_0_0_wdata(ram_w8_l4096_id0_0_0_wdata),
    .ram_w8_l4096_id0_0_0_wenable(ram_w8_l4096_id0_0_0_wenable),
    .ram_w8_l4096_id0_0_0_enable(ram_w8_l4096_id0_0_0_enable),
    .ram_w8_l4096_id0_0_1_addr(ram_w8_l4096_id0_0_1_addr),
    .ram_w8_l4096_id0_0_1_rdata(ram_w8_l4096_id0_0_1_rdata),
    .ram_w8_l4096_id0_0_1_wdata(ram_w8_l4096_id0_0_1_wdata),
    .ram_w8_l4096_id0_0_1_wenable(ram_w8_l4096_id0_0_1_wenable),
    .ram_w8_l4096_id0_0_1_enable(ram_w8_l4096_id0_0_1_enable)
  );

  wire [10-1:0] ram_w8_l4096_id0_1_0_addr;
  wire [8-1:0] ram_w8_l4096_id0_1_0_rdata;
  wire [8-1:0] ram_w8_l4096_id0_1_0_wdata;
  wire ram_w8_l4096_id0_1_0_wenable;
  wire ram_w8_l4096_id0_1_0_enable;
  wire [10-1:0] ram_w8_l4096_id0_1_1_addr;
  wire [8-1:0] ram_w8_l4096_id0_1_1_rdata;
  wire [8-1:0] ram_w8_l4096_id0_1_1_wdata;
  wire ram_w8_l4096_id0_1_1_wenable;
  wire ram_w8_l4096_id0_1_1_enable;
  assign ram_w8_l4096_id0_1_0_wdata = 'hx;
  assign ram_w8_l4096_id0_1_0_wenable = 0;

  ram_w8_l4096_id0_1
  inst_ram_w8_l4096_id0_1
  (
    .CLK(CLK),
    .ram_w8_l4096_id0_1_0_addr(ram_w8_l4096_id0_1_0_addr),
    .ram_w8_l4096_id0_1_0_rdata(ram_w8_l4096_id0_1_0_rdata),
    .ram_w8_l4096_id0_1_0_wdata(ram_w8_l4096_id0_1_0_wdata),
    .ram_w8_l4096_id0_1_0_wenable(ram_w8_l4096_id0_1_0_wenable),
    .ram_w8_l4096_id0_1_0_enable(ram_w8_l4096_id0_1_0_enable),
    .ram_w8_l4096_id0_1_1_addr(ram_w8_l4096_id0_1_1_addr),
    .ram_w8_l4096_id0_1_1_rdata(ram_w8_l4096_id0_1_1_rdata),
    .ram_w8_l4096_id0_1_1_wdata(ram_w8_l4096_id0_1_1_wdata),
    .ram_w8_l4096_id0_1_1_wenable(ram_w8_l4096_id0_1_1_wenable),
    .ram_w8_l4096_id0_1_1_enable(ram_w8_l4096_id0_1_1_enable)
  );

  wire [10-1:0] ram_w8_l4096_id0_2_0_addr;
  wire [8-1:0] ram_w8_l4096_id0_2_0_rdata;
  wire [8-1:0] ram_w8_l4096_id0_2_0_wdata;
  wire ram_w8_l4096_id0_2_0_wenable;
  wire ram_w8_l4096_id0_2_0_enable;
  wire [10-1:0] ram_w8_l4096_id0_2_1_addr;
  wire [8-1:0] ram_w8_l4096_id0_2_1_rdata;
  wire [8-1:0] ram_w8_l4096_id0_2_1_wdata;
  wire ram_w8_l4096_id0_2_1_wenable;
  wire ram_w8_l4096_id0_2_1_enable;
  assign ram_w8_l4096_id0_2_0_wdata = 'hx;
  assign ram_w8_l4096_id0_2_0_wenable = 0;

  ram_w8_l4096_id0_2
  inst_ram_w8_l4096_id0_2
  (
    .CLK(CLK),
    .ram_w8_l4096_id0_2_0_addr(ram_w8_l4096_id0_2_0_addr),
    .ram_w8_l4096_id0_2_0_rdata(ram_w8_l4096_id0_2_0_rdata),
    .ram_w8_l4096_id0_2_0_wdata(ram_w8_l4096_id0_2_0_wdata),
    .ram_w8_l4096_id0_2_0_wenable(ram_w8_l4096_id0_2_0_wenable),
    .ram_w8_l4096_id0_2_0_enable(ram_w8_l4096_id0_2_0_enable),
    .ram_w8_l4096_id0_2_1_addr(ram_w8_l4096_id0_2_1_addr),
    .ram_w8_l4096_id0_2_1_rdata(ram_w8_l4096_id0_2_1_rdata),
    .ram_w8_l4096_id0_2_1_wdata(ram_w8_l4096_id0_2_1_wdata),
    .ram_w8_l4096_id0_2_1_wenable(ram_w8_l4096_id0_2_1_wenable),
    .ram_w8_l4096_id0_2_1_enable(ram_w8_l4096_id0_2_1_enable)
  );

  wire [10-1:0] ram_w8_l4096_id0_3_0_addr;
  wire [8-1:0] ram_w8_l4096_id0_3_0_rdata;
  wire [8-1:0] ram_w8_l4096_id0_3_0_wdata;
  wire ram_w8_l4096_id0_3_0_wenable;
  wire ram_w8_l4096_id0_3_0_enable;
  wire [10-1:0] ram_w8_l4096_id0_3_1_addr;
  wire [8-1:0] ram_w8_l4096_id0_3_1_rdata;
  wire [8-1:0] ram_w8_l4096_id0_3_1_wdata;
  wire ram_w8_l4096_id0_3_1_wenable;
  wire ram_w8_l4096_id0_3_1_enable;
  assign ram_w8_l4096_id0_3_0_wdata = 'hx;
  assign ram_w8_l4096_id0_3_0_wenable = 0;

  ram_w8_l4096_id0_3
  inst_ram_w8_l4096_id0_3
  (
    .CLK(CLK),
    .ram_w8_l4096_id0_3_0_addr(ram_w8_l4096_id0_3_0_addr),
    .ram_w8_l4096_id0_3_0_rdata(ram_w8_l4096_id0_3_0_rdata),
    .ram_w8_l4096_id0_3_0_wdata(ram_w8_l4096_id0_3_0_wdata),
    .ram_w8_l4096_id0_3_0_wenable(ram_w8_l4096_id0_3_0_wenable),
    .ram_w8_l4096_id0_3_0_enable(ram_w8_l4096_id0_3_0_enable),
    .ram_w8_l4096_id0_3_1_addr(ram_w8_l4096_id0_3_1_addr),
    .ram_w8_l4096_id0_3_1_rdata(ram_w8_l4096_id0_3_1_rdata),
    .ram_w8_l4096_id0_3_1_wdata(ram_w8_l4096_id0_3_1_wdata),
    .ram_w8_l4096_id0_3_1_wenable(ram_w8_l4096_id0_3_1_wenable),
    .ram_w8_l4096_id0_3_1_enable(ram_w8_l4096_id0_3_1_enable)
  );

  wire [10-1:0] ram_w8_l4096_id1_0_0_addr;
  wire [8-1:0] ram_w8_l4096_id1_0_0_rdata;
  wire [8-1:0] ram_w8_l4096_id1_0_0_wdata;
  wire ram_w8_l4096_id1_0_0_wenable;
  wire ram_w8_l4096_id1_0_0_enable;
  wire [10-1:0] ram_w8_l4096_id1_0_1_addr;
  wire [8-1:0] ram_w8_l4096_id1_0_1_rdata;
  wire [8-1:0] ram_w8_l4096_id1_0_1_wdata;
  wire ram_w8_l4096_id1_0_1_wenable;
  wire ram_w8_l4096_id1_0_1_enable;
  assign ram_w8_l4096_id1_0_0_wdata = 'hx;
  assign ram_w8_l4096_id1_0_0_wenable = 0;

  ram_w8_l4096_id1_0
  inst_ram_w8_l4096_id1_0
  (
    .CLK(CLK),
    .ram_w8_l4096_id1_0_0_addr(ram_w8_l4096_id1_0_0_addr),
    .ram_w8_l4096_id1_0_0_rdata(ram_w8_l4096_id1_0_0_rdata),
    .ram_w8_l4096_id1_0_0_wdata(ram_w8_l4096_id1_0_0_wdata),
    .ram_w8_l4096_id1_0_0_wenable(ram_w8_l4096_id1_0_0_wenable),
    .ram_w8_l4096_id1_0_0_enable(ram_w8_l4096_id1_0_0_enable),
    .ram_w8_l4096_id1_0_1_addr(ram_w8_l4096_id1_0_1_addr),
    .ram_w8_l4096_id1_0_1_rdata(ram_w8_l4096_id1_0_1_rdata),
    .ram_w8_l4096_id1_0_1_wdata(ram_w8_l4096_id1_0_1_wdata),
    .ram_w8_l4096_id1_0_1_wenable(ram_w8_l4096_id1_0_1_wenable),
    .ram_w8_l4096_id1_0_1_enable(ram_w8_l4096_id1_0_1_enable)
  );

  wire [10-1:0] ram_w8_l4096_id1_1_0_addr;
  wire [8-1:0] ram_w8_l4096_id1_1_0_rdata;
  wire [8-1:0] ram_w8_l4096_id1_1_0_wdata;
  wire ram_w8_l4096_id1_1_0_wenable;
  wire ram_w8_l4096_id1_1_0_enable;
  wire [10-1:0] ram_w8_l4096_id1_1_1_addr;
  wire [8-1:0] ram_w8_l4096_id1_1_1_rdata;
  wire [8-1:0] ram_w8_l4096_id1_1_1_wdata;
  wire ram_w8_l4096_id1_1_1_wenable;
  wire ram_w8_l4096_id1_1_1_enable;
  assign ram_w8_l4096_id1_1_0_wdata = 'hx;
  assign ram_w8_l4096_id1_1_0_wenable = 0;

  ram_w8_l4096_id1_1
  inst_ram_w8_l4096_id1_1
  (
    .CLK(CLK),
    .ram_w8_l4096_id1_1_0_addr(ram_w8_l4096_id1_1_0_addr),
    .ram_w8_l4096_id1_1_0_rdata(ram_w8_l4096_id1_1_0_rdata),
    .ram_w8_l4096_id1_1_0_wdata(ram_w8_l4096_id1_1_0_wdata),
    .ram_w8_l4096_id1_1_0_wenable(ram_w8_l4096_id1_1_0_wenable),
    .ram_w8_l4096_id1_1_0_enable(ram_w8_l4096_id1_1_0_enable),
    .ram_w8_l4096_id1_1_1_addr(ram_w8_l4096_id1_1_1_addr),
    .ram_w8_l4096_id1_1_1_rdata(ram_w8_l4096_id1_1_1_rdata),
    .ram_w8_l4096_id1_1_1_wdata(ram_w8_l4096_id1_1_1_wdata),
    .ram_w8_l4096_id1_1_1_wenable(ram_w8_l4096_id1_1_1_wenable),
    .ram_w8_l4096_id1_1_1_enable(ram_w8_l4096_id1_1_1_enable)
  );

  wire [10-1:0] ram_w8_l4096_id1_2_0_addr;
  wire [8-1:0] ram_w8_l4096_id1_2_0_rdata;
  wire [8-1:0] ram_w8_l4096_id1_2_0_wdata;
  wire ram_w8_l4096_id1_2_0_wenable;
  wire ram_w8_l4096_id1_2_0_enable;
  wire [10-1:0] ram_w8_l4096_id1_2_1_addr;
  wire [8-1:0] ram_w8_l4096_id1_2_1_rdata;
  wire [8-1:0] ram_w8_l4096_id1_2_1_wdata;
  wire ram_w8_l4096_id1_2_1_wenable;
  wire ram_w8_l4096_id1_2_1_enable;
  assign ram_w8_l4096_id1_2_0_wdata = 'hx;
  assign ram_w8_l4096_id1_2_0_wenable = 0;

  ram_w8_l4096_id1_2
  inst_ram_w8_l4096_id1_2
  (
    .CLK(CLK),
    .ram_w8_l4096_id1_2_0_addr(ram_w8_l4096_id1_2_0_addr),
    .ram_w8_l4096_id1_2_0_rdata(ram_w8_l4096_id1_2_0_rdata),
    .ram_w8_l4096_id1_2_0_wdata(ram_w8_l4096_id1_2_0_wdata),
    .ram_w8_l4096_id1_2_0_wenable(ram_w8_l4096_id1_2_0_wenable),
    .ram_w8_l4096_id1_2_0_enable(ram_w8_l4096_id1_2_0_enable),
    .ram_w8_l4096_id1_2_1_addr(ram_w8_l4096_id1_2_1_addr),
    .ram_w8_l4096_id1_2_1_rdata(ram_w8_l4096_id1_2_1_rdata),
    .ram_w8_l4096_id1_2_1_wdata(ram_w8_l4096_id1_2_1_wdata),
    .ram_w8_l4096_id1_2_1_wenable(ram_w8_l4096_id1_2_1_wenable),
    .ram_w8_l4096_id1_2_1_enable(ram_w8_l4096_id1_2_1_enable)
  );

  wire [10-1:0] ram_w8_l4096_id1_3_0_addr;
  wire [8-1:0] ram_w8_l4096_id1_3_0_rdata;
  wire [8-1:0] ram_w8_l4096_id1_3_0_wdata;
  wire ram_w8_l4096_id1_3_0_wenable;
  wire ram_w8_l4096_id1_3_0_enable;
  wire [10-1:0] ram_w8_l4096_id1_3_1_addr;
  wire [8-1:0] ram_w8_l4096_id1_3_1_rdata;
  wire [8-1:0] ram_w8_l4096_id1_3_1_wdata;
  wire ram_w8_l4096_id1_3_1_wenable;
  wire ram_w8_l4096_id1_3_1_enable;
  assign ram_w8_l4096_id1_3_0_wdata = 'hx;
  assign ram_w8_l4096_id1_3_0_wenable = 0;

  ram_w8_l4096_id1_3
  inst_ram_w8_l4096_id1_3
  (
    .CLK(CLK),
    .ram_w8_l4096_id1_3_0_addr(ram_w8_l4096_id1_3_0_addr),
    .ram_w8_l4096_id1_3_0_rdata(ram_w8_l4096_id1_3_0_rdata),
    .ram_w8_l4096_id1_3_0_wdata(ram_w8_l4096_id1_3_0_wdata),
    .ram_w8_l4096_id1_3_0_wenable(ram_w8_l4096_id1_3_0_wenable),
    .ram_w8_l4096_id1_3_0_enable(ram_w8_l4096_id1_3_0_enable),
    .ram_w8_l4096_id1_3_1_addr(ram_w8_l4096_id1_3_1_addr),
    .ram_w8_l4096_id1_3_1_rdata(ram_w8_l4096_id1_3_1_rdata),
    .ram_w8_l4096_id1_3_1_wdata(ram_w8_l4096_id1_3_1_wdata),
    .ram_w8_l4096_id1_3_1_wenable(ram_w8_l4096_id1_3_1_wenable),
    .ram_w8_l4096_id1_3_1_enable(ram_w8_l4096_id1_3_1_enable)
  );

  wire [10-1:0] ram_w8_l4096_id2_0_0_addr;
  wire [8-1:0] ram_w8_l4096_id2_0_0_rdata;
  wire [8-1:0] ram_w8_l4096_id2_0_0_wdata;
  wire ram_w8_l4096_id2_0_0_wenable;
  wire ram_w8_l4096_id2_0_0_enable;
  wire [10-1:0] ram_w8_l4096_id2_0_1_addr;
  wire [8-1:0] ram_w8_l4096_id2_0_1_rdata;
  wire [8-1:0] ram_w8_l4096_id2_0_1_wdata;
  wire ram_w8_l4096_id2_0_1_wenable;
  wire ram_w8_l4096_id2_0_1_enable;
  assign ram_w8_l4096_id2_0_0_wdata = 'hx;
  assign ram_w8_l4096_id2_0_0_wenable = 0;

  ram_w8_l4096_id2_0
  inst_ram_w8_l4096_id2_0
  (
    .CLK(CLK),
    .ram_w8_l4096_id2_0_0_addr(ram_w8_l4096_id2_0_0_addr),
    .ram_w8_l4096_id2_0_0_rdata(ram_w8_l4096_id2_0_0_rdata),
    .ram_w8_l4096_id2_0_0_wdata(ram_w8_l4096_id2_0_0_wdata),
    .ram_w8_l4096_id2_0_0_wenable(ram_w8_l4096_id2_0_0_wenable),
    .ram_w8_l4096_id2_0_0_enable(ram_w8_l4096_id2_0_0_enable),
    .ram_w8_l4096_id2_0_1_addr(ram_w8_l4096_id2_0_1_addr),
    .ram_w8_l4096_id2_0_1_rdata(ram_w8_l4096_id2_0_1_rdata),
    .ram_w8_l4096_id2_0_1_wdata(ram_w8_l4096_id2_0_1_wdata),
    .ram_w8_l4096_id2_0_1_wenable(ram_w8_l4096_id2_0_1_wenable),
    .ram_w8_l4096_id2_0_1_enable(ram_w8_l4096_id2_0_1_enable)
  );

  wire [10-1:0] ram_w8_l4096_id2_1_0_addr;
  wire [8-1:0] ram_w8_l4096_id2_1_0_rdata;
  wire [8-1:0] ram_w8_l4096_id2_1_0_wdata;
  wire ram_w8_l4096_id2_1_0_wenable;
  wire ram_w8_l4096_id2_1_0_enable;
  wire [10-1:0] ram_w8_l4096_id2_1_1_addr;
  wire [8-1:0] ram_w8_l4096_id2_1_1_rdata;
  wire [8-1:0] ram_w8_l4096_id2_1_1_wdata;
  wire ram_w8_l4096_id2_1_1_wenable;
  wire ram_w8_l4096_id2_1_1_enable;
  assign ram_w8_l4096_id2_1_0_wdata = 'hx;
  assign ram_w8_l4096_id2_1_0_wenable = 0;

  ram_w8_l4096_id2_1
  inst_ram_w8_l4096_id2_1
  (
    .CLK(CLK),
    .ram_w8_l4096_id2_1_0_addr(ram_w8_l4096_id2_1_0_addr),
    .ram_w8_l4096_id2_1_0_rdata(ram_w8_l4096_id2_1_0_rdata),
    .ram_w8_l4096_id2_1_0_wdata(ram_w8_l4096_id2_1_0_wdata),
    .ram_w8_l4096_id2_1_0_wenable(ram_w8_l4096_id2_1_0_wenable),
    .ram_w8_l4096_id2_1_0_enable(ram_w8_l4096_id2_1_0_enable),
    .ram_w8_l4096_id2_1_1_addr(ram_w8_l4096_id2_1_1_addr),
    .ram_w8_l4096_id2_1_1_rdata(ram_w8_l4096_id2_1_1_rdata),
    .ram_w8_l4096_id2_1_1_wdata(ram_w8_l4096_id2_1_1_wdata),
    .ram_w8_l4096_id2_1_1_wenable(ram_w8_l4096_id2_1_1_wenable),
    .ram_w8_l4096_id2_1_1_enable(ram_w8_l4096_id2_1_1_enable)
  );

  wire [10-1:0] ram_w8_l4096_id2_2_0_addr;
  wire [8-1:0] ram_w8_l4096_id2_2_0_rdata;
  wire [8-1:0] ram_w8_l4096_id2_2_0_wdata;
  wire ram_w8_l4096_id2_2_0_wenable;
  wire ram_w8_l4096_id2_2_0_enable;
  wire [10-1:0] ram_w8_l4096_id2_2_1_addr;
  wire [8-1:0] ram_w8_l4096_id2_2_1_rdata;
  wire [8-1:0] ram_w8_l4096_id2_2_1_wdata;
  wire ram_w8_l4096_id2_2_1_wenable;
  wire ram_w8_l4096_id2_2_1_enable;
  assign ram_w8_l4096_id2_2_0_wdata = 'hx;
  assign ram_w8_l4096_id2_2_0_wenable = 0;

  ram_w8_l4096_id2_2
  inst_ram_w8_l4096_id2_2
  (
    .CLK(CLK),
    .ram_w8_l4096_id2_2_0_addr(ram_w8_l4096_id2_2_0_addr),
    .ram_w8_l4096_id2_2_0_rdata(ram_w8_l4096_id2_2_0_rdata),
    .ram_w8_l4096_id2_2_0_wdata(ram_w8_l4096_id2_2_0_wdata),
    .ram_w8_l4096_id2_2_0_wenable(ram_w8_l4096_id2_2_0_wenable),
    .ram_w8_l4096_id2_2_0_enable(ram_w8_l4096_id2_2_0_enable),
    .ram_w8_l4096_id2_2_1_addr(ram_w8_l4096_id2_2_1_addr),
    .ram_w8_l4096_id2_2_1_rdata(ram_w8_l4096_id2_2_1_rdata),
    .ram_w8_l4096_id2_2_1_wdata(ram_w8_l4096_id2_2_1_wdata),
    .ram_w8_l4096_id2_2_1_wenable(ram_w8_l4096_id2_2_1_wenable),
    .ram_w8_l4096_id2_2_1_enable(ram_w8_l4096_id2_2_1_enable)
  );

  wire [10-1:0] ram_w8_l4096_id2_3_0_addr;
  wire [8-1:0] ram_w8_l4096_id2_3_0_rdata;
  wire [8-1:0] ram_w8_l4096_id2_3_0_wdata;
  wire ram_w8_l4096_id2_3_0_wenable;
  wire ram_w8_l4096_id2_3_0_enable;
  wire [10-1:0] ram_w8_l4096_id2_3_1_addr;
  wire [8-1:0] ram_w8_l4096_id2_3_1_rdata;
  wire [8-1:0] ram_w8_l4096_id2_3_1_wdata;
  wire ram_w8_l4096_id2_3_1_wenable;
  wire ram_w8_l4096_id2_3_1_enable;
  assign ram_w8_l4096_id2_3_0_wdata = 'hx;
  assign ram_w8_l4096_id2_3_0_wenable = 0;

  ram_w8_l4096_id2_3
  inst_ram_w8_l4096_id2_3
  (
    .CLK(CLK),
    .ram_w8_l4096_id2_3_0_addr(ram_w8_l4096_id2_3_0_addr),
    .ram_w8_l4096_id2_3_0_rdata(ram_w8_l4096_id2_3_0_rdata),
    .ram_w8_l4096_id2_3_0_wdata(ram_w8_l4096_id2_3_0_wdata),
    .ram_w8_l4096_id2_3_0_wenable(ram_w8_l4096_id2_3_0_wenable),
    .ram_w8_l4096_id2_3_0_enable(ram_w8_l4096_id2_3_0_enable),
    .ram_w8_l4096_id2_3_1_addr(ram_w8_l4096_id2_3_1_addr),
    .ram_w8_l4096_id2_3_1_rdata(ram_w8_l4096_id2_3_1_rdata),
    .ram_w8_l4096_id2_3_1_wdata(ram_w8_l4096_id2_3_1_wdata),
    .ram_w8_l4096_id2_3_1_wenable(ram_w8_l4096_id2_3_1_wenable),
    .ram_w8_l4096_id2_3_1_enable(ram_w8_l4096_id2_3_1_enable)
  );

  wire [10-1:0] ram_w8_l4096_id3_0_0_addr;
  wire [8-1:0] ram_w8_l4096_id3_0_0_rdata;
  wire [8-1:0] ram_w8_l4096_id3_0_0_wdata;
  wire ram_w8_l4096_id3_0_0_wenable;
  wire ram_w8_l4096_id3_0_0_enable;
  wire [10-1:0] ram_w8_l4096_id3_0_1_addr;
  wire [8-1:0] ram_w8_l4096_id3_0_1_rdata;
  wire [8-1:0] ram_w8_l4096_id3_0_1_wdata;
  wire ram_w8_l4096_id3_0_1_wenable;
  wire ram_w8_l4096_id3_0_1_enable;
  assign ram_w8_l4096_id3_0_0_wdata = 'hx;
  assign ram_w8_l4096_id3_0_0_wenable = 0;

  ram_w8_l4096_id3_0
  inst_ram_w8_l4096_id3_0
  (
    .CLK(CLK),
    .ram_w8_l4096_id3_0_0_addr(ram_w8_l4096_id3_0_0_addr),
    .ram_w8_l4096_id3_0_0_rdata(ram_w8_l4096_id3_0_0_rdata),
    .ram_w8_l4096_id3_0_0_wdata(ram_w8_l4096_id3_0_0_wdata),
    .ram_w8_l4096_id3_0_0_wenable(ram_w8_l4096_id3_0_0_wenable),
    .ram_w8_l4096_id3_0_0_enable(ram_w8_l4096_id3_0_0_enable),
    .ram_w8_l4096_id3_0_1_addr(ram_w8_l4096_id3_0_1_addr),
    .ram_w8_l4096_id3_0_1_rdata(ram_w8_l4096_id3_0_1_rdata),
    .ram_w8_l4096_id3_0_1_wdata(ram_w8_l4096_id3_0_1_wdata),
    .ram_w8_l4096_id3_0_1_wenable(ram_w8_l4096_id3_0_1_wenable),
    .ram_w8_l4096_id3_0_1_enable(ram_w8_l4096_id3_0_1_enable)
  );

  wire [10-1:0] ram_w8_l4096_id3_1_0_addr;
  wire [8-1:0] ram_w8_l4096_id3_1_0_rdata;
  wire [8-1:0] ram_w8_l4096_id3_1_0_wdata;
  wire ram_w8_l4096_id3_1_0_wenable;
  wire ram_w8_l4096_id3_1_0_enable;
  wire [10-1:0] ram_w8_l4096_id3_1_1_addr;
  wire [8-1:0] ram_w8_l4096_id3_1_1_rdata;
  wire [8-1:0] ram_w8_l4096_id3_1_1_wdata;
  wire ram_w8_l4096_id3_1_1_wenable;
  wire ram_w8_l4096_id3_1_1_enable;
  assign ram_w8_l4096_id3_1_0_wdata = 'hx;
  assign ram_w8_l4096_id3_1_0_wenable = 0;

  ram_w8_l4096_id3_1
  inst_ram_w8_l4096_id3_1
  (
    .CLK(CLK),
    .ram_w8_l4096_id3_1_0_addr(ram_w8_l4096_id3_1_0_addr),
    .ram_w8_l4096_id3_1_0_rdata(ram_w8_l4096_id3_1_0_rdata),
    .ram_w8_l4096_id3_1_0_wdata(ram_w8_l4096_id3_1_0_wdata),
    .ram_w8_l4096_id3_1_0_wenable(ram_w8_l4096_id3_1_0_wenable),
    .ram_w8_l4096_id3_1_0_enable(ram_w8_l4096_id3_1_0_enable),
    .ram_w8_l4096_id3_1_1_addr(ram_w8_l4096_id3_1_1_addr),
    .ram_w8_l4096_id3_1_1_rdata(ram_w8_l4096_id3_1_1_rdata),
    .ram_w8_l4096_id3_1_1_wdata(ram_w8_l4096_id3_1_1_wdata),
    .ram_w8_l4096_id3_1_1_wenable(ram_w8_l4096_id3_1_1_wenable),
    .ram_w8_l4096_id3_1_1_enable(ram_w8_l4096_id3_1_1_enable)
  );

  wire [10-1:0] ram_w8_l4096_id3_2_0_addr;
  wire [8-1:0] ram_w8_l4096_id3_2_0_rdata;
  wire [8-1:0] ram_w8_l4096_id3_2_0_wdata;
  wire ram_w8_l4096_id3_2_0_wenable;
  wire ram_w8_l4096_id3_2_0_enable;
  wire [10-1:0] ram_w8_l4096_id3_2_1_addr;
  wire [8-1:0] ram_w8_l4096_id3_2_1_rdata;
  wire [8-1:0] ram_w8_l4096_id3_2_1_wdata;
  wire ram_w8_l4096_id3_2_1_wenable;
  wire ram_w8_l4096_id3_2_1_enable;
  assign ram_w8_l4096_id3_2_0_wdata = 'hx;
  assign ram_w8_l4096_id3_2_0_wenable = 0;

  ram_w8_l4096_id3_2
  inst_ram_w8_l4096_id3_2
  (
    .CLK(CLK),
    .ram_w8_l4096_id3_2_0_addr(ram_w8_l4096_id3_2_0_addr),
    .ram_w8_l4096_id3_2_0_rdata(ram_w8_l4096_id3_2_0_rdata),
    .ram_w8_l4096_id3_2_0_wdata(ram_w8_l4096_id3_2_0_wdata),
    .ram_w8_l4096_id3_2_0_wenable(ram_w8_l4096_id3_2_0_wenable),
    .ram_w8_l4096_id3_2_0_enable(ram_w8_l4096_id3_2_0_enable),
    .ram_w8_l4096_id3_2_1_addr(ram_w8_l4096_id3_2_1_addr),
    .ram_w8_l4096_id3_2_1_rdata(ram_w8_l4096_id3_2_1_rdata),
    .ram_w8_l4096_id3_2_1_wdata(ram_w8_l4096_id3_2_1_wdata),
    .ram_w8_l4096_id3_2_1_wenable(ram_w8_l4096_id3_2_1_wenable),
    .ram_w8_l4096_id3_2_1_enable(ram_w8_l4096_id3_2_1_enable)
  );

  wire [10-1:0] ram_w8_l4096_id3_3_0_addr;
  wire [8-1:0] ram_w8_l4096_id3_3_0_rdata;
  wire [8-1:0] ram_w8_l4096_id3_3_0_wdata;
  wire ram_w8_l4096_id3_3_0_wenable;
  wire ram_w8_l4096_id3_3_0_enable;
  wire [10-1:0] ram_w8_l4096_id3_3_1_addr;
  wire [8-1:0] ram_w8_l4096_id3_3_1_rdata;
  wire [8-1:0] ram_w8_l4096_id3_3_1_wdata;
  wire ram_w8_l4096_id3_3_1_wenable;
  wire ram_w8_l4096_id3_3_1_enable;
  assign ram_w8_l4096_id3_3_0_wdata = 'hx;
  assign ram_w8_l4096_id3_3_0_wenable = 0;

  ram_w8_l4096_id3_3
  inst_ram_w8_l4096_id3_3
  (
    .CLK(CLK),
    .ram_w8_l4096_id3_3_0_addr(ram_w8_l4096_id3_3_0_addr),
    .ram_w8_l4096_id3_3_0_rdata(ram_w8_l4096_id3_3_0_rdata),
    .ram_w8_l4096_id3_3_0_wdata(ram_w8_l4096_id3_3_0_wdata),
    .ram_w8_l4096_id3_3_0_wenable(ram_w8_l4096_id3_3_0_wenable),
    .ram_w8_l4096_id3_3_0_enable(ram_w8_l4096_id3_3_0_enable),
    .ram_w8_l4096_id3_3_1_addr(ram_w8_l4096_id3_3_1_addr),
    .ram_w8_l4096_id3_3_1_rdata(ram_w8_l4096_id3_3_1_rdata),
    .ram_w8_l4096_id3_3_1_wdata(ram_w8_l4096_id3_3_1_wdata),
    .ram_w8_l4096_id3_3_1_wenable(ram_w8_l4096_id3_3_1_wenable),
    .ram_w8_l4096_id3_3_1_enable(ram_w8_l4096_id3_3_1_enable)
  );

  wire [10-1:0] ram_w8_l4096_id4_0_0_addr;
  wire [8-1:0] ram_w8_l4096_id4_0_0_rdata;
  wire [8-1:0] ram_w8_l4096_id4_0_0_wdata;
  wire ram_w8_l4096_id4_0_0_wenable;
  wire ram_w8_l4096_id4_0_0_enable;
  wire [10-1:0] ram_w8_l4096_id4_0_1_addr;
  wire [8-1:0] ram_w8_l4096_id4_0_1_rdata;
  wire [8-1:0] ram_w8_l4096_id4_0_1_wdata;
  wire ram_w8_l4096_id4_0_1_wenable;
  wire ram_w8_l4096_id4_0_1_enable;
  assign ram_w8_l4096_id4_0_0_wdata = 'hx;
  assign ram_w8_l4096_id4_0_0_wenable = 0;

  ram_w8_l4096_id4_0
  inst_ram_w8_l4096_id4_0
  (
    .CLK(CLK),
    .ram_w8_l4096_id4_0_0_addr(ram_w8_l4096_id4_0_0_addr),
    .ram_w8_l4096_id4_0_0_rdata(ram_w8_l4096_id4_0_0_rdata),
    .ram_w8_l4096_id4_0_0_wdata(ram_w8_l4096_id4_0_0_wdata),
    .ram_w8_l4096_id4_0_0_wenable(ram_w8_l4096_id4_0_0_wenable),
    .ram_w8_l4096_id4_0_0_enable(ram_w8_l4096_id4_0_0_enable),
    .ram_w8_l4096_id4_0_1_addr(ram_w8_l4096_id4_0_1_addr),
    .ram_w8_l4096_id4_0_1_rdata(ram_w8_l4096_id4_0_1_rdata),
    .ram_w8_l4096_id4_0_1_wdata(ram_w8_l4096_id4_0_1_wdata),
    .ram_w8_l4096_id4_0_1_wenable(ram_w8_l4096_id4_0_1_wenable),
    .ram_w8_l4096_id4_0_1_enable(ram_w8_l4096_id4_0_1_enable)
  );

  wire [10-1:0] ram_w8_l4096_id4_1_0_addr;
  wire [8-1:0] ram_w8_l4096_id4_1_0_rdata;
  wire [8-1:0] ram_w8_l4096_id4_1_0_wdata;
  wire ram_w8_l4096_id4_1_0_wenable;
  wire ram_w8_l4096_id4_1_0_enable;
  wire [10-1:0] ram_w8_l4096_id4_1_1_addr;
  wire [8-1:0] ram_w8_l4096_id4_1_1_rdata;
  wire [8-1:0] ram_w8_l4096_id4_1_1_wdata;
  wire ram_w8_l4096_id4_1_1_wenable;
  wire ram_w8_l4096_id4_1_1_enable;
  assign ram_w8_l4096_id4_1_0_wdata = 'hx;
  assign ram_w8_l4096_id4_1_0_wenable = 0;

  ram_w8_l4096_id4_1
  inst_ram_w8_l4096_id4_1
  (
    .CLK(CLK),
    .ram_w8_l4096_id4_1_0_addr(ram_w8_l4096_id4_1_0_addr),
    .ram_w8_l4096_id4_1_0_rdata(ram_w8_l4096_id4_1_0_rdata),
    .ram_w8_l4096_id4_1_0_wdata(ram_w8_l4096_id4_1_0_wdata),
    .ram_w8_l4096_id4_1_0_wenable(ram_w8_l4096_id4_1_0_wenable),
    .ram_w8_l4096_id4_1_0_enable(ram_w8_l4096_id4_1_0_enable),
    .ram_w8_l4096_id4_1_1_addr(ram_w8_l4096_id4_1_1_addr),
    .ram_w8_l4096_id4_1_1_rdata(ram_w8_l4096_id4_1_1_rdata),
    .ram_w8_l4096_id4_1_1_wdata(ram_w8_l4096_id4_1_1_wdata),
    .ram_w8_l4096_id4_1_1_wenable(ram_w8_l4096_id4_1_1_wenable),
    .ram_w8_l4096_id4_1_1_enable(ram_w8_l4096_id4_1_1_enable)
  );

  wire [10-1:0] ram_w8_l4096_id4_2_0_addr;
  wire [8-1:0] ram_w8_l4096_id4_2_0_rdata;
  wire [8-1:0] ram_w8_l4096_id4_2_0_wdata;
  wire ram_w8_l4096_id4_2_0_wenable;
  wire ram_w8_l4096_id4_2_0_enable;
  wire [10-1:0] ram_w8_l4096_id4_2_1_addr;
  wire [8-1:0] ram_w8_l4096_id4_2_1_rdata;
  wire [8-1:0] ram_w8_l4096_id4_2_1_wdata;
  wire ram_w8_l4096_id4_2_1_wenable;
  wire ram_w8_l4096_id4_2_1_enable;
  assign ram_w8_l4096_id4_2_0_wdata = 'hx;
  assign ram_w8_l4096_id4_2_0_wenable = 0;

  ram_w8_l4096_id4_2
  inst_ram_w8_l4096_id4_2
  (
    .CLK(CLK),
    .ram_w8_l4096_id4_2_0_addr(ram_w8_l4096_id4_2_0_addr),
    .ram_w8_l4096_id4_2_0_rdata(ram_w8_l4096_id4_2_0_rdata),
    .ram_w8_l4096_id4_2_0_wdata(ram_w8_l4096_id4_2_0_wdata),
    .ram_w8_l4096_id4_2_0_wenable(ram_w8_l4096_id4_2_0_wenable),
    .ram_w8_l4096_id4_2_0_enable(ram_w8_l4096_id4_2_0_enable),
    .ram_w8_l4096_id4_2_1_addr(ram_w8_l4096_id4_2_1_addr),
    .ram_w8_l4096_id4_2_1_rdata(ram_w8_l4096_id4_2_1_rdata),
    .ram_w8_l4096_id4_2_1_wdata(ram_w8_l4096_id4_2_1_wdata),
    .ram_w8_l4096_id4_2_1_wenable(ram_w8_l4096_id4_2_1_wenable),
    .ram_w8_l4096_id4_2_1_enable(ram_w8_l4096_id4_2_1_enable)
  );

  wire [10-1:0] ram_w8_l4096_id4_3_0_addr;
  wire [8-1:0] ram_w8_l4096_id4_3_0_rdata;
  wire [8-1:0] ram_w8_l4096_id4_3_0_wdata;
  wire ram_w8_l4096_id4_3_0_wenable;
  wire ram_w8_l4096_id4_3_0_enable;
  wire [10-1:0] ram_w8_l4096_id4_3_1_addr;
  wire [8-1:0] ram_w8_l4096_id4_3_1_rdata;
  wire [8-1:0] ram_w8_l4096_id4_3_1_wdata;
  wire ram_w8_l4096_id4_3_1_wenable;
  wire ram_w8_l4096_id4_3_1_enable;
  assign ram_w8_l4096_id4_3_0_wdata = 'hx;
  assign ram_w8_l4096_id4_3_0_wenable = 0;

  ram_w8_l4096_id4_3
  inst_ram_w8_l4096_id4_3
  (
    .CLK(CLK),
    .ram_w8_l4096_id4_3_0_addr(ram_w8_l4096_id4_3_0_addr),
    .ram_w8_l4096_id4_3_0_rdata(ram_w8_l4096_id4_3_0_rdata),
    .ram_w8_l4096_id4_3_0_wdata(ram_w8_l4096_id4_3_0_wdata),
    .ram_w8_l4096_id4_3_0_wenable(ram_w8_l4096_id4_3_0_wenable),
    .ram_w8_l4096_id4_3_0_enable(ram_w8_l4096_id4_3_0_enable),
    .ram_w8_l4096_id4_3_1_addr(ram_w8_l4096_id4_3_1_addr),
    .ram_w8_l4096_id4_3_1_rdata(ram_w8_l4096_id4_3_1_rdata),
    .ram_w8_l4096_id4_3_1_wdata(ram_w8_l4096_id4_3_1_wdata),
    .ram_w8_l4096_id4_3_1_wenable(ram_w8_l4096_id4_3_1_wenable),
    .ram_w8_l4096_id4_3_1_enable(ram_w8_l4096_id4_3_1_enable)
  );

  wire [10-1:0] ram_w8_l4096_id5_0_0_addr;
  wire [8-1:0] ram_w8_l4096_id5_0_0_rdata;
  wire [8-1:0] ram_w8_l4096_id5_0_0_wdata;
  wire ram_w8_l4096_id5_0_0_wenable;
  wire ram_w8_l4096_id5_0_0_enable;
  wire [10-1:0] ram_w8_l4096_id5_0_1_addr;
  wire [8-1:0] ram_w8_l4096_id5_0_1_rdata;
  wire [8-1:0] ram_w8_l4096_id5_0_1_wdata;
  wire ram_w8_l4096_id5_0_1_wenable;
  wire ram_w8_l4096_id5_0_1_enable;
  assign ram_w8_l4096_id5_0_0_wdata = 'hx;
  assign ram_w8_l4096_id5_0_0_wenable = 0;

  ram_w8_l4096_id5_0
  inst_ram_w8_l4096_id5_0
  (
    .CLK(CLK),
    .ram_w8_l4096_id5_0_0_addr(ram_w8_l4096_id5_0_0_addr),
    .ram_w8_l4096_id5_0_0_rdata(ram_w8_l4096_id5_0_0_rdata),
    .ram_w8_l4096_id5_0_0_wdata(ram_w8_l4096_id5_0_0_wdata),
    .ram_w8_l4096_id5_0_0_wenable(ram_w8_l4096_id5_0_0_wenable),
    .ram_w8_l4096_id5_0_0_enable(ram_w8_l4096_id5_0_0_enable),
    .ram_w8_l4096_id5_0_1_addr(ram_w8_l4096_id5_0_1_addr),
    .ram_w8_l4096_id5_0_1_rdata(ram_w8_l4096_id5_0_1_rdata),
    .ram_w8_l4096_id5_0_1_wdata(ram_w8_l4096_id5_0_1_wdata),
    .ram_w8_l4096_id5_0_1_wenable(ram_w8_l4096_id5_0_1_wenable),
    .ram_w8_l4096_id5_0_1_enable(ram_w8_l4096_id5_0_1_enable)
  );

  wire [10-1:0] ram_w8_l4096_id5_1_0_addr;
  wire [8-1:0] ram_w8_l4096_id5_1_0_rdata;
  wire [8-1:0] ram_w8_l4096_id5_1_0_wdata;
  wire ram_w8_l4096_id5_1_0_wenable;
  wire ram_w8_l4096_id5_1_0_enable;
  wire [10-1:0] ram_w8_l4096_id5_1_1_addr;
  wire [8-1:0] ram_w8_l4096_id5_1_1_rdata;
  wire [8-1:0] ram_w8_l4096_id5_1_1_wdata;
  wire ram_w8_l4096_id5_1_1_wenable;
  wire ram_w8_l4096_id5_1_1_enable;
  assign ram_w8_l4096_id5_1_0_wdata = 'hx;
  assign ram_w8_l4096_id5_1_0_wenable = 0;

  ram_w8_l4096_id5_1
  inst_ram_w8_l4096_id5_1
  (
    .CLK(CLK),
    .ram_w8_l4096_id5_1_0_addr(ram_w8_l4096_id5_1_0_addr),
    .ram_w8_l4096_id5_1_0_rdata(ram_w8_l4096_id5_1_0_rdata),
    .ram_w8_l4096_id5_1_0_wdata(ram_w8_l4096_id5_1_0_wdata),
    .ram_w8_l4096_id5_1_0_wenable(ram_w8_l4096_id5_1_0_wenable),
    .ram_w8_l4096_id5_1_0_enable(ram_w8_l4096_id5_1_0_enable),
    .ram_w8_l4096_id5_1_1_addr(ram_w8_l4096_id5_1_1_addr),
    .ram_w8_l4096_id5_1_1_rdata(ram_w8_l4096_id5_1_1_rdata),
    .ram_w8_l4096_id5_1_1_wdata(ram_w8_l4096_id5_1_1_wdata),
    .ram_w8_l4096_id5_1_1_wenable(ram_w8_l4096_id5_1_1_wenable),
    .ram_w8_l4096_id5_1_1_enable(ram_w8_l4096_id5_1_1_enable)
  );

  wire [10-1:0] ram_w8_l4096_id5_2_0_addr;
  wire [8-1:0] ram_w8_l4096_id5_2_0_rdata;
  wire [8-1:0] ram_w8_l4096_id5_2_0_wdata;
  wire ram_w8_l4096_id5_2_0_wenable;
  wire ram_w8_l4096_id5_2_0_enable;
  wire [10-1:0] ram_w8_l4096_id5_2_1_addr;
  wire [8-1:0] ram_w8_l4096_id5_2_1_rdata;
  wire [8-1:0] ram_w8_l4096_id5_2_1_wdata;
  wire ram_w8_l4096_id5_2_1_wenable;
  wire ram_w8_l4096_id5_2_1_enable;
  assign ram_w8_l4096_id5_2_0_wdata = 'hx;
  assign ram_w8_l4096_id5_2_0_wenable = 0;

  ram_w8_l4096_id5_2
  inst_ram_w8_l4096_id5_2
  (
    .CLK(CLK),
    .ram_w8_l4096_id5_2_0_addr(ram_w8_l4096_id5_2_0_addr),
    .ram_w8_l4096_id5_2_0_rdata(ram_w8_l4096_id5_2_0_rdata),
    .ram_w8_l4096_id5_2_0_wdata(ram_w8_l4096_id5_2_0_wdata),
    .ram_w8_l4096_id5_2_0_wenable(ram_w8_l4096_id5_2_0_wenable),
    .ram_w8_l4096_id5_2_0_enable(ram_w8_l4096_id5_2_0_enable),
    .ram_w8_l4096_id5_2_1_addr(ram_w8_l4096_id5_2_1_addr),
    .ram_w8_l4096_id5_2_1_rdata(ram_w8_l4096_id5_2_1_rdata),
    .ram_w8_l4096_id5_2_1_wdata(ram_w8_l4096_id5_2_1_wdata),
    .ram_w8_l4096_id5_2_1_wenable(ram_w8_l4096_id5_2_1_wenable),
    .ram_w8_l4096_id5_2_1_enable(ram_w8_l4096_id5_2_1_enable)
  );

  wire [10-1:0] ram_w8_l4096_id5_3_0_addr;
  wire [8-1:0] ram_w8_l4096_id5_3_0_rdata;
  wire [8-1:0] ram_w8_l4096_id5_3_0_wdata;
  wire ram_w8_l4096_id5_3_0_wenable;
  wire ram_w8_l4096_id5_3_0_enable;
  wire [10-1:0] ram_w8_l4096_id5_3_1_addr;
  wire [8-1:0] ram_w8_l4096_id5_3_1_rdata;
  wire [8-1:0] ram_w8_l4096_id5_3_1_wdata;
  wire ram_w8_l4096_id5_3_1_wenable;
  wire ram_w8_l4096_id5_3_1_enable;
  assign ram_w8_l4096_id5_3_0_wdata = 'hx;
  assign ram_w8_l4096_id5_3_0_wenable = 0;

  ram_w8_l4096_id5_3
  inst_ram_w8_l4096_id5_3
  (
    .CLK(CLK),
    .ram_w8_l4096_id5_3_0_addr(ram_w8_l4096_id5_3_0_addr),
    .ram_w8_l4096_id5_3_0_rdata(ram_w8_l4096_id5_3_0_rdata),
    .ram_w8_l4096_id5_3_0_wdata(ram_w8_l4096_id5_3_0_wdata),
    .ram_w8_l4096_id5_3_0_wenable(ram_w8_l4096_id5_3_0_wenable),
    .ram_w8_l4096_id5_3_0_enable(ram_w8_l4096_id5_3_0_enable),
    .ram_w8_l4096_id5_3_1_addr(ram_w8_l4096_id5_3_1_addr),
    .ram_w8_l4096_id5_3_1_rdata(ram_w8_l4096_id5_3_1_rdata),
    .ram_w8_l4096_id5_3_1_wdata(ram_w8_l4096_id5_3_1_wdata),
    .ram_w8_l4096_id5_3_1_wenable(ram_w8_l4096_id5_3_1_wenable),
    .ram_w8_l4096_id5_3_1_enable(ram_w8_l4096_id5_3_1_enable)
  );

  wire [10-1:0] ram_w8_l4096_id6_0_0_addr;
  wire [8-1:0] ram_w8_l4096_id6_0_0_rdata;
  wire [8-1:0] ram_w8_l4096_id6_0_0_wdata;
  wire ram_w8_l4096_id6_0_0_wenable;
  wire ram_w8_l4096_id6_0_0_enable;
  wire [10-1:0] ram_w8_l4096_id6_0_1_addr;
  wire [8-1:0] ram_w8_l4096_id6_0_1_rdata;
  wire [8-1:0] ram_w8_l4096_id6_0_1_wdata;
  wire ram_w8_l4096_id6_0_1_wenable;
  wire ram_w8_l4096_id6_0_1_enable;
  assign ram_w8_l4096_id6_0_0_wdata = 'hx;
  assign ram_w8_l4096_id6_0_0_wenable = 0;

  ram_w8_l4096_id6_0
  inst_ram_w8_l4096_id6_0
  (
    .CLK(CLK),
    .ram_w8_l4096_id6_0_0_addr(ram_w8_l4096_id6_0_0_addr),
    .ram_w8_l4096_id6_0_0_rdata(ram_w8_l4096_id6_0_0_rdata),
    .ram_w8_l4096_id6_0_0_wdata(ram_w8_l4096_id6_0_0_wdata),
    .ram_w8_l4096_id6_0_0_wenable(ram_w8_l4096_id6_0_0_wenable),
    .ram_w8_l4096_id6_0_0_enable(ram_w8_l4096_id6_0_0_enable),
    .ram_w8_l4096_id6_0_1_addr(ram_w8_l4096_id6_0_1_addr),
    .ram_w8_l4096_id6_0_1_rdata(ram_w8_l4096_id6_0_1_rdata),
    .ram_w8_l4096_id6_0_1_wdata(ram_w8_l4096_id6_0_1_wdata),
    .ram_w8_l4096_id6_0_1_wenable(ram_w8_l4096_id6_0_1_wenable),
    .ram_w8_l4096_id6_0_1_enable(ram_w8_l4096_id6_0_1_enable)
  );

  wire [10-1:0] ram_w8_l4096_id6_1_0_addr;
  wire [8-1:0] ram_w8_l4096_id6_1_0_rdata;
  wire [8-1:0] ram_w8_l4096_id6_1_0_wdata;
  wire ram_w8_l4096_id6_1_0_wenable;
  wire ram_w8_l4096_id6_1_0_enable;
  wire [10-1:0] ram_w8_l4096_id6_1_1_addr;
  wire [8-1:0] ram_w8_l4096_id6_1_1_rdata;
  wire [8-1:0] ram_w8_l4096_id6_1_1_wdata;
  wire ram_w8_l4096_id6_1_1_wenable;
  wire ram_w8_l4096_id6_1_1_enable;
  assign ram_w8_l4096_id6_1_0_wdata = 'hx;
  assign ram_w8_l4096_id6_1_0_wenable = 0;

  ram_w8_l4096_id6_1
  inst_ram_w8_l4096_id6_1
  (
    .CLK(CLK),
    .ram_w8_l4096_id6_1_0_addr(ram_w8_l4096_id6_1_0_addr),
    .ram_w8_l4096_id6_1_0_rdata(ram_w8_l4096_id6_1_0_rdata),
    .ram_w8_l4096_id6_1_0_wdata(ram_w8_l4096_id6_1_0_wdata),
    .ram_w8_l4096_id6_1_0_wenable(ram_w8_l4096_id6_1_0_wenable),
    .ram_w8_l4096_id6_1_0_enable(ram_w8_l4096_id6_1_0_enable),
    .ram_w8_l4096_id6_1_1_addr(ram_w8_l4096_id6_1_1_addr),
    .ram_w8_l4096_id6_1_1_rdata(ram_w8_l4096_id6_1_1_rdata),
    .ram_w8_l4096_id6_1_1_wdata(ram_w8_l4096_id6_1_1_wdata),
    .ram_w8_l4096_id6_1_1_wenable(ram_w8_l4096_id6_1_1_wenable),
    .ram_w8_l4096_id6_1_1_enable(ram_w8_l4096_id6_1_1_enable)
  );

  wire [10-1:0] ram_w8_l4096_id6_2_0_addr;
  wire [8-1:0] ram_w8_l4096_id6_2_0_rdata;
  wire [8-1:0] ram_w8_l4096_id6_2_0_wdata;
  wire ram_w8_l4096_id6_2_0_wenable;
  wire ram_w8_l4096_id6_2_0_enable;
  wire [10-1:0] ram_w8_l4096_id6_2_1_addr;
  wire [8-1:0] ram_w8_l4096_id6_2_1_rdata;
  wire [8-1:0] ram_w8_l4096_id6_2_1_wdata;
  wire ram_w8_l4096_id6_2_1_wenable;
  wire ram_w8_l4096_id6_2_1_enable;
  assign ram_w8_l4096_id6_2_0_wdata = 'hx;
  assign ram_w8_l4096_id6_2_0_wenable = 0;

  ram_w8_l4096_id6_2
  inst_ram_w8_l4096_id6_2
  (
    .CLK(CLK),
    .ram_w8_l4096_id6_2_0_addr(ram_w8_l4096_id6_2_0_addr),
    .ram_w8_l4096_id6_2_0_rdata(ram_w8_l4096_id6_2_0_rdata),
    .ram_w8_l4096_id6_2_0_wdata(ram_w8_l4096_id6_2_0_wdata),
    .ram_w8_l4096_id6_2_0_wenable(ram_w8_l4096_id6_2_0_wenable),
    .ram_w8_l4096_id6_2_0_enable(ram_w8_l4096_id6_2_0_enable),
    .ram_w8_l4096_id6_2_1_addr(ram_w8_l4096_id6_2_1_addr),
    .ram_w8_l4096_id6_2_1_rdata(ram_w8_l4096_id6_2_1_rdata),
    .ram_w8_l4096_id6_2_1_wdata(ram_w8_l4096_id6_2_1_wdata),
    .ram_w8_l4096_id6_2_1_wenable(ram_w8_l4096_id6_2_1_wenable),
    .ram_w8_l4096_id6_2_1_enable(ram_w8_l4096_id6_2_1_enable)
  );

  wire [10-1:0] ram_w8_l4096_id6_3_0_addr;
  wire [8-1:0] ram_w8_l4096_id6_3_0_rdata;
  wire [8-1:0] ram_w8_l4096_id6_3_0_wdata;
  wire ram_w8_l4096_id6_3_0_wenable;
  wire ram_w8_l4096_id6_3_0_enable;
  wire [10-1:0] ram_w8_l4096_id6_3_1_addr;
  wire [8-1:0] ram_w8_l4096_id6_3_1_rdata;
  wire [8-1:0] ram_w8_l4096_id6_3_1_wdata;
  wire ram_w8_l4096_id6_3_1_wenable;
  wire ram_w8_l4096_id6_3_1_enable;
  assign ram_w8_l4096_id6_3_0_wdata = 'hx;
  assign ram_w8_l4096_id6_3_0_wenable = 0;

  ram_w8_l4096_id6_3
  inst_ram_w8_l4096_id6_3
  (
    .CLK(CLK),
    .ram_w8_l4096_id6_3_0_addr(ram_w8_l4096_id6_3_0_addr),
    .ram_w8_l4096_id6_3_0_rdata(ram_w8_l4096_id6_3_0_rdata),
    .ram_w8_l4096_id6_3_0_wdata(ram_w8_l4096_id6_3_0_wdata),
    .ram_w8_l4096_id6_3_0_wenable(ram_w8_l4096_id6_3_0_wenable),
    .ram_w8_l4096_id6_3_0_enable(ram_w8_l4096_id6_3_0_enable),
    .ram_w8_l4096_id6_3_1_addr(ram_w8_l4096_id6_3_1_addr),
    .ram_w8_l4096_id6_3_1_rdata(ram_w8_l4096_id6_3_1_rdata),
    .ram_w8_l4096_id6_3_1_wdata(ram_w8_l4096_id6_3_1_wdata),
    .ram_w8_l4096_id6_3_1_wenable(ram_w8_l4096_id6_3_1_wenable),
    .ram_w8_l4096_id6_3_1_enable(ram_w8_l4096_id6_3_1_enable)
  );

  wire [10-1:0] ram_w8_l4096_id7_0_0_addr;
  wire [8-1:0] ram_w8_l4096_id7_0_0_rdata;
  wire [8-1:0] ram_w8_l4096_id7_0_0_wdata;
  wire ram_w8_l4096_id7_0_0_wenable;
  wire ram_w8_l4096_id7_0_0_enable;
  wire [10-1:0] ram_w8_l4096_id7_0_1_addr;
  wire [8-1:0] ram_w8_l4096_id7_0_1_rdata;
  wire [8-1:0] ram_w8_l4096_id7_0_1_wdata;
  wire ram_w8_l4096_id7_0_1_wenable;
  wire ram_w8_l4096_id7_0_1_enable;
  assign ram_w8_l4096_id7_0_0_wdata = 'hx;
  assign ram_w8_l4096_id7_0_0_wenable = 0;

  ram_w8_l4096_id7_0
  inst_ram_w8_l4096_id7_0
  (
    .CLK(CLK),
    .ram_w8_l4096_id7_0_0_addr(ram_w8_l4096_id7_0_0_addr),
    .ram_w8_l4096_id7_0_0_rdata(ram_w8_l4096_id7_0_0_rdata),
    .ram_w8_l4096_id7_0_0_wdata(ram_w8_l4096_id7_0_0_wdata),
    .ram_w8_l4096_id7_0_0_wenable(ram_w8_l4096_id7_0_0_wenable),
    .ram_w8_l4096_id7_0_0_enable(ram_w8_l4096_id7_0_0_enable),
    .ram_w8_l4096_id7_0_1_addr(ram_w8_l4096_id7_0_1_addr),
    .ram_w8_l4096_id7_0_1_rdata(ram_w8_l4096_id7_0_1_rdata),
    .ram_w8_l4096_id7_0_1_wdata(ram_w8_l4096_id7_0_1_wdata),
    .ram_w8_l4096_id7_0_1_wenable(ram_w8_l4096_id7_0_1_wenable),
    .ram_w8_l4096_id7_0_1_enable(ram_w8_l4096_id7_0_1_enable)
  );

  wire [10-1:0] ram_w8_l4096_id7_1_0_addr;
  wire [8-1:0] ram_w8_l4096_id7_1_0_rdata;
  wire [8-1:0] ram_w8_l4096_id7_1_0_wdata;
  wire ram_w8_l4096_id7_1_0_wenable;
  wire ram_w8_l4096_id7_1_0_enable;
  wire [10-1:0] ram_w8_l4096_id7_1_1_addr;
  wire [8-1:0] ram_w8_l4096_id7_1_1_rdata;
  wire [8-1:0] ram_w8_l4096_id7_1_1_wdata;
  wire ram_w8_l4096_id7_1_1_wenable;
  wire ram_w8_l4096_id7_1_1_enable;
  assign ram_w8_l4096_id7_1_0_wdata = 'hx;
  assign ram_w8_l4096_id7_1_0_wenable = 0;

  ram_w8_l4096_id7_1
  inst_ram_w8_l4096_id7_1
  (
    .CLK(CLK),
    .ram_w8_l4096_id7_1_0_addr(ram_w8_l4096_id7_1_0_addr),
    .ram_w8_l4096_id7_1_0_rdata(ram_w8_l4096_id7_1_0_rdata),
    .ram_w8_l4096_id7_1_0_wdata(ram_w8_l4096_id7_1_0_wdata),
    .ram_w8_l4096_id7_1_0_wenable(ram_w8_l4096_id7_1_0_wenable),
    .ram_w8_l4096_id7_1_0_enable(ram_w8_l4096_id7_1_0_enable),
    .ram_w8_l4096_id7_1_1_addr(ram_w8_l4096_id7_1_1_addr),
    .ram_w8_l4096_id7_1_1_rdata(ram_w8_l4096_id7_1_1_rdata),
    .ram_w8_l4096_id7_1_1_wdata(ram_w8_l4096_id7_1_1_wdata),
    .ram_w8_l4096_id7_1_1_wenable(ram_w8_l4096_id7_1_1_wenable),
    .ram_w8_l4096_id7_1_1_enable(ram_w8_l4096_id7_1_1_enable)
  );

  wire [10-1:0] ram_w8_l4096_id7_2_0_addr;
  wire [8-1:0] ram_w8_l4096_id7_2_0_rdata;
  wire [8-1:0] ram_w8_l4096_id7_2_0_wdata;
  wire ram_w8_l4096_id7_2_0_wenable;
  wire ram_w8_l4096_id7_2_0_enable;
  wire [10-1:0] ram_w8_l4096_id7_2_1_addr;
  wire [8-1:0] ram_w8_l4096_id7_2_1_rdata;
  wire [8-1:0] ram_w8_l4096_id7_2_1_wdata;
  wire ram_w8_l4096_id7_2_1_wenable;
  wire ram_w8_l4096_id7_2_1_enable;
  assign ram_w8_l4096_id7_2_0_wdata = 'hx;
  assign ram_w8_l4096_id7_2_0_wenable = 0;

  ram_w8_l4096_id7_2
  inst_ram_w8_l4096_id7_2
  (
    .CLK(CLK),
    .ram_w8_l4096_id7_2_0_addr(ram_w8_l4096_id7_2_0_addr),
    .ram_w8_l4096_id7_2_0_rdata(ram_w8_l4096_id7_2_0_rdata),
    .ram_w8_l4096_id7_2_0_wdata(ram_w8_l4096_id7_2_0_wdata),
    .ram_w8_l4096_id7_2_0_wenable(ram_w8_l4096_id7_2_0_wenable),
    .ram_w8_l4096_id7_2_0_enable(ram_w8_l4096_id7_2_0_enable),
    .ram_w8_l4096_id7_2_1_addr(ram_w8_l4096_id7_2_1_addr),
    .ram_w8_l4096_id7_2_1_rdata(ram_w8_l4096_id7_2_1_rdata),
    .ram_w8_l4096_id7_2_1_wdata(ram_w8_l4096_id7_2_1_wdata),
    .ram_w8_l4096_id7_2_1_wenable(ram_w8_l4096_id7_2_1_wenable),
    .ram_w8_l4096_id7_2_1_enable(ram_w8_l4096_id7_2_1_enable)
  );

  wire [10-1:0] ram_w8_l4096_id7_3_0_addr;
  wire [8-1:0] ram_w8_l4096_id7_3_0_rdata;
  wire [8-1:0] ram_w8_l4096_id7_3_0_wdata;
  wire ram_w8_l4096_id7_3_0_wenable;
  wire ram_w8_l4096_id7_3_0_enable;
  wire [10-1:0] ram_w8_l4096_id7_3_1_addr;
  wire [8-1:0] ram_w8_l4096_id7_3_1_rdata;
  wire [8-1:0] ram_w8_l4096_id7_3_1_wdata;
  wire ram_w8_l4096_id7_3_1_wenable;
  wire ram_w8_l4096_id7_3_1_enable;
  assign ram_w8_l4096_id7_3_0_wdata = 'hx;
  assign ram_w8_l4096_id7_3_0_wenable = 0;

  ram_w8_l4096_id7_3
  inst_ram_w8_l4096_id7_3
  (
    .CLK(CLK),
    .ram_w8_l4096_id7_3_0_addr(ram_w8_l4096_id7_3_0_addr),
    .ram_w8_l4096_id7_3_0_rdata(ram_w8_l4096_id7_3_0_rdata),
    .ram_w8_l4096_id7_3_0_wdata(ram_w8_l4096_id7_3_0_wdata),
    .ram_w8_l4096_id7_3_0_wenable(ram_w8_l4096_id7_3_0_wenable),
    .ram_w8_l4096_id7_3_0_enable(ram_w8_l4096_id7_3_0_enable),
    .ram_w8_l4096_id7_3_1_addr(ram_w8_l4096_id7_3_1_addr),
    .ram_w8_l4096_id7_3_1_rdata(ram_w8_l4096_id7_3_1_rdata),
    .ram_w8_l4096_id7_3_1_wdata(ram_w8_l4096_id7_3_1_wdata),
    .ram_w8_l4096_id7_3_1_wenable(ram_w8_l4096_id7_3_1_wenable),
    .ram_w8_l4096_id7_3_1_enable(ram_w8_l4096_id7_3_1_enable)
  );

  wire [10-1:0] ram_w8_l4096_id8_0_0_addr;
  wire [8-1:0] ram_w8_l4096_id8_0_0_rdata;
  wire [8-1:0] ram_w8_l4096_id8_0_0_wdata;
  wire ram_w8_l4096_id8_0_0_wenable;
  wire ram_w8_l4096_id8_0_0_enable;
  wire [10-1:0] ram_w8_l4096_id8_0_1_addr;
  wire [8-1:0] ram_w8_l4096_id8_0_1_rdata;
  wire [8-1:0] ram_w8_l4096_id8_0_1_wdata;
  wire ram_w8_l4096_id8_0_1_wenable;
  wire ram_w8_l4096_id8_0_1_enable;
  assign ram_w8_l4096_id8_0_0_wdata = 'hx;
  assign ram_w8_l4096_id8_0_0_wenable = 0;

  ram_w8_l4096_id8_0
  inst_ram_w8_l4096_id8_0
  (
    .CLK(CLK),
    .ram_w8_l4096_id8_0_0_addr(ram_w8_l4096_id8_0_0_addr),
    .ram_w8_l4096_id8_0_0_rdata(ram_w8_l4096_id8_0_0_rdata),
    .ram_w8_l4096_id8_0_0_wdata(ram_w8_l4096_id8_0_0_wdata),
    .ram_w8_l4096_id8_0_0_wenable(ram_w8_l4096_id8_0_0_wenable),
    .ram_w8_l4096_id8_0_0_enable(ram_w8_l4096_id8_0_0_enable),
    .ram_w8_l4096_id8_0_1_addr(ram_w8_l4096_id8_0_1_addr),
    .ram_w8_l4096_id8_0_1_rdata(ram_w8_l4096_id8_0_1_rdata),
    .ram_w8_l4096_id8_0_1_wdata(ram_w8_l4096_id8_0_1_wdata),
    .ram_w8_l4096_id8_0_1_wenable(ram_w8_l4096_id8_0_1_wenable),
    .ram_w8_l4096_id8_0_1_enable(ram_w8_l4096_id8_0_1_enable)
  );

  wire [10-1:0] ram_w8_l4096_id8_1_0_addr;
  wire [8-1:0] ram_w8_l4096_id8_1_0_rdata;
  wire [8-1:0] ram_w8_l4096_id8_1_0_wdata;
  wire ram_w8_l4096_id8_1_0_wenable;
  wire ram_w8_l4096_id8_1_0_enable;
  wire [10-1:0] ram_w8_l4096_id8_1_1_addr;
  wire [8-1:0] ram_w8_l4096_id8_1_1_rdata;
  wire [8-1:0] ram_w8_l4096_id8_1_1_wdata;
  wire ram_w8_l4096_id8_1_1_wenable;
  wire ram_w8_l4096_id8_1_1_enable;
  assign ram_w8_l4096_id8_1_0_wdata = 'hx;
  assign ram_w8_l4096_id8_1_0_wenable = 0;

  ram_w8_l4096_id8_1
  inst_ram_w8_l4096_id8_1
  (
    .CLK(CLK),
    .ram_w8_l4096_id8_1_0_addr(ram_w8_l4096_id8_1_0_addr),
    .ram_w8_l4096_id8_1_0_rdata(ram_w8_l4096_id8_1_0_rdata),
    .ram_w8_l4096_id8_1_0_wdata(ram_w8_l4096_id8_1_0_wdata),
    .ram_w8_l4096_id8_1_0_wenable(ram_w8_l4096_id8_1_0_wenable),
    .ram_w8_l4096_id8_1_0_enable(ram_w8_l4096_id8_1_0_enable),
    .ram_w8_l4096_id8_1_1_addr(ram_w8_l4096_id8_1_1_addr),
    .ram_w8_l4096_id8_1_1_rdata(ram_w8_l4096_id8_1_1_rdata),
    .ram_w8_l4096_id8_1_1_wdata(ram_w8_l4096_id8_1_1_wdata),
    .ram_w8_l4096_id8_1_1_wenable(ram_w8_l4096_id8_1_1_wenable),
    .ram_w8_l4096_id8_1_1_enable(ram_w8_l4096_id8_1_1_enable)
  );

  wire [10-1:0] ram_w8_l4096_id8_2_0_addr;
  wire [8-1:0] ram_w8_l4096_id8_2_0_rdata;
  wire [8-1:0] ram_w8_l4096_id8_2_0_wdata;
  wire ram_w8_l4096_id8_2_0_wenable;
  wire ram_w8_l4096_id8_2_0_enable;
  wire [10-1:0] ram_w8_l4096_id8_2_1_addr;
  wire [8-1:0] ram_w8_l4096_id8_2_1_rdata;
  wire [8-1:0] ram_w8_l4096_id8_2_1_wdata;
  wire ram_w8_l4096_id8_2_1_wenable;
  wire ram_w8_l4096_id8_2_1_enable;
  assign ram_w8_l4096_id8_2_0_wdata = 'hx;
  assign ram_w8_l4096_id8_2_0_wenable = 0;

  ram_w8_l4096_id8_2
  inst_ram_w8_l4096_id8_2
  (
    .CLK(CLK),
    .ram_w8_l4096_id8_2_0_addr(ram_w8_l4096_id8_2_0_addr),
    .ram_w8_l4096_id8_2_0_rdata(ram_w8_l4096_id8_2_0_rdata),
    .ram_w8_l4096_id8_2_0_wdata(ram_w8_l4096_id8_2_0_wdata),
    .ram_w8_l4096_id8_2_0_wenable(ram_w8_l4096_id8_2_0_wenable),
    .ram_w8_l4096_id8_2_0_enable(ram_w8_l4096_id8_2_0_enable),
    .ram_w8_l4096_id8_2_1_addr(ram_w8_l4096_id8_2_1_addr),
    .ram_w8_l4096_id8_2_1_rdata(ram_w8_l4096_id8_2_1_rdata),
    .ram_w8_l4096_id8_2_1_wdata(ram_w8_l4096_id8_2_1_wdata),
    .ram_w8_l4096_id8_2_1_wenable(ram_w8_l4096_id8_2_1_wenable),
    .ram_w8_l4096_id8_2_1_enable(ram_w8_l4096_id8_2_1_enable)
  );

  wire [10-1:0] ram_w8_l4096_id8_3_0_addr;
  wire [8-1:0] ram_w8_l4096_id8_3_0_rdata;
  wire [8-1:0] ram_w8_l4096_id8_3_0_wdata;
  wire ram_w8_l4096_id8_3_0_wenable;
  wire ram_w8_l4096_id8_3_0_enable;
  wire [10-1:0] ram_w8_l4096_id8_3_1_addr;
  wire [8-1:0] ram_w8_l4096_id8_3_1_rdata;
  wire [8-1:0] ram_w8_l4096_id8_3_1_wdata;
  wire ram_w8_l4096_id8_3_1_wenable;
  wire ram_w8_l4096_id8_3_1_enable;
  assign ram_w8_l4096_id8_3_0_wdata = 'hx;
  assign ram_w8_l4096_id8_3_0_wenable = 0;

  ram_w8_l4096_id8_3
  inst_ram_w8_l4096_id8_3
  (
    .CLK(CLK),
    .ram_w8_l4096_id8_3_0_addr(ram_w8_l4096_id8_3_0_addr),
    .ram_w8_l4096_id8_3_0_rdata(ram_w8_l4096_id8_3_0_rdata),
    .ram_w8_l4096_id8_3_0_wdata(ram_w8_l4096_id8_3_0_wdata),
    .ram_w8_l4096_id8_3_0_wenable(ram_w8_l4096_id8_3_0_wenable),
    .ram_w8_l4096_id8_3_0_enable(ram_w8_l4096_id8_3_0_enable),
    .ram_w8_l4096_id8_3_1_addr(ram_w8_l4096_id8_3_1_addr),
    .ram_w8_l4096_id8_3_1_rdata(ram_w8_l4096_id8_3_1_rdata),
    .ram_w8_l4096_id8_3_1_wdata(ram_w8_l4096_id8_3_1_wdata),
    .ram_w8_l4096_id8_3_1_wenable(ram_w8_l4096_id8_3_1_wenable),
    .ram_w8_l4096_id8_3_1_enable(ram_w8_l4096_id8_3_1_enable)
  );

  wire [9-1:0] ram_w8_l2048_id0_0_0_addr;
  wire [8-1:0] ram_w8_l2048_id0_0_0_rdata;
  wire [8-1:0] ram_w8_l2048_id0_0_0_wdata;
  wire ram_w8_l2048_id0_0_0_wenable;
  wire ram_w8_l2048_id0_0_0_enable;
  wire [9-1:0] ram_w8_l2048_id0_0_1_addr;
  wire [8-1:0] ram_w8_l2048_id0_0_1_rdata;
  wire [8-1:0] ram_w8_l2048_id0_0_1_wdata;
  wire ram_w8_l2048_id0_0_1_wenable;
  wire ram_w8_l2048_id0_0_1_enable;
  assign ram_w8_l2048_id0_0_0_wdata = 'hx;
  assign ram_w8_l2048_id0_0_0_wenable = 0;

  ram_w8_l2048_id0_0
  inst_ram_w8_l2048_id0_0
  (
    .CLK(CLK),
    .ram_w8_l2048_id0_0_0_addr(ram_w8_l2048_id0_0_0_addr),
    .ram_w8_l2048_id0_0_0_rdata(ram_w8_l2048_id0_0_0_rdata),
    .ram_w8_l2048_id0_0_0_wdata(ram_w8_l2048_id0_0_0_wdata),
    .ram_w8_l2048_id0_0_0_wenable(ram_w8_l2048_id0_0_0_wenable),
    .ram_w8_l2048_id0_0_0_enable(ram_w8_l2048_id0_0_0_enable),
    .ram_w8_l2048_id0_0_1_addr(ram_w8_l2048_id0_0_1_addr),
    .ram_w8_l2048_id0_0_1_rdata(ram_w8_l2048_id0_0_1_rdata),
    .ram_w8_l2048_id0_0_1_wdata(ram_w8_l2048_id0_0_1_wdata),
    .ram_w8_l2048_id0_0_1_wenable(ram_w8_l2048_id0_0_1_wenable),
    .ram_w8_l2048_id0_0_1_enable(ram_w8_l2048_id0_0_1_enable)
  );

  wire [9-1:0] ram_w8_l2048_id0_1_0_addr;
  wire [8-1:0] ram_w8_l2048_id0_1_0_rdata;
  wire [8-1:0] ram_w8_l2048_id0_1_0_wdata;
  wire ram_w8_l2048_id0_1_0_wenable;
  wire ram_w8_l2048_id0_1_0_enable;
  wire [9-1:0] ram_w8_l2048_id0_1_1_addr;
  wire [8-1:0] ram_w8_l2048_id0_1_1_rdata;
  wire [8-1:0] ram_w8_l2048_id0_1_1_wdata;
  wire ram_w8_l2048_id0_1_1_wenable;
  wire ram_w8_l2048_id0_1_1_enable;
  assign ram_w8_l2048_id0_1_0_wdata = 'hx;
  assign ram_w8_l2048_id0_1_0_wenable = 0;

  ram_w8_l2048_id0_1
  inst_ram_w8_l2048_id0_1
  (
    .CLK(CLK),
    .ram_w8_l2048_id0_1_0_addr(ram_w8_l2048_id0_1_0_addr),
    .ram_w8_l2048_id0_1_0_rdata(ram_w8_l2048_id0_1_0_rdata),
    .ram_w8_l2048_id0_1_0_wdata(ram_w8_l2048_id0_1_0_wdata),
    .ram_w8_l2048_id0_1_0_wenable(ram_w8_l2048_id0_1_0_wenable),
    .ram_w8_l2048_id0_1_0_enable(ram_w8_l2048_id0_1_0_enable),
    .ram_w8_l2048_id0_1_1_addr(ram_w8_l2048_id0_1_1_addr),
    .ram_w8_l2048_id0_1_1_rdata(ram_w8_l2048_id0_1_1_rdata),
    .ram_w8_l2048_id0_1_1_wdata(ram_w8_l2048_id0_1_1_wdata),
    .ram_w8_l2048_id0_1_1_wenable(ram_w8_l2048_id0_1_1_wenable),
    .ram_w8_l2048_id0_1_1_enable(ram_w8_l2048_id0_1_1_enable)
  );

  wire [9-1:0] ram_w8_l2048_id0_2_0_addr;
  wire [8-1:0] ram_w8_l2048_id0_2_0_rdata;
  wire [8-1:0] ram_w8_l2048_id0_2_0_wdata;
  wire ram_w8_l2048_id0_2_0_wenable;
  wire ram_w8_l2048_id0_2_0_enable;
  wire [9-1:0] ram_w8_l2048_id0_2_1_addr;
  wire [8-1:0] ram_w8_l2048_id0_2_1_rdata;
  wire [8-1:0] ram_w8_l2048_id0_2_1_wdata;
  wire ram_w8_l2048_id0_2_1_wenable;
  wire ram_w8_l2048_id0_2_1_enable;
  assign ram_w8_l2048_id0_2_0_wdata = 'hx;
  assign ram_w8_l2048_id0_2_0_wenable = 0;

  ram_w8_l2048_id0_2
  inst_ram_w8_l2048_id0_2
  (
    .CLK(CLK),
    .ram_w8_l2048_id0_2_0_addr(ram_w8_l2048_id0_2_0_addr),
    .ram_w8_l2048_id0_2_0_rdata(ram_w8_l2048_id0_2_0_rdata),
    .ram_w8_l2048_id0_2_0_wdata(ram_w8_l2048_id0_2_0_wdata),
    .ram_w8_l2048_id0_2_0_wenable(ram_w8_l2048_id0_2_0_wenable),
    .ram_w8_l2048_id0_2_0_enable(ram_w8_l2048_id0_2_0_enable),
    .ram_w8_l2048_id0_2_1_addr(ram_w8_l2048_id0_2_1_addr),
    .ram_w8_l2048_id0_2_1_rdata(ram_w8_l2048_id0_2_1_rdata),
    .ram_w8_l2048_id0_2_1_wdata(ram_w8_l2048_id0_2_1_wdata),
    .ram_w8_l2048_id0_2_1_wenable(ram_w8_l2048_id0_2_1_wenable),
    .ram_w8_l2048_id0_2_1_enable(ram_w8_l2048_id0_2_1_enable)
  );

  wire [9-1:0] ram_w8_l2048_id0_3_0_addr;
  wire [8-1:0] ram_w8_l2048_id0_3_0_rdata;
  wire [8-1:0] ram_w8_l2048_id0_3_0_wdata;
  wire ram_w8_l2048_id0_3_0_wenable;
  wire ram_w8_l2048_id0_3_0_enable;
  wire [9-1:0] ram_w8_l2048_id0_3_1_addr;
  wire [8-1:0] ram_w8_l2048_id0_3_1_rdata;
  wire [8-1:0] ram_w8_l2048_id0_3_1_wdata;
  wire ram_w8_l2048_id0_3_1_wenable;
  wire ram_w8_l2048_id0_3_1_enable;
  assign ram_w8_l2048_id0_3_0_wdata = 'hx;
  assign ram_w8_l2048_id0_3_0_wenable = 0;

  ram_w8_l2048_id0_3
  inst_ram_w8_l2048_id0_3
  (
    .CLK(CLK),
    .ram_w8_l2048_id0_3_0_addr(ram_w8_l2048_id0_3_0_addr),
    .ram_w8_l2048_id0_3_0_rdata(ram_w8_l2048_id0_3_0_rdata),
    .ram_w8_l2048_id0_3_0_wdata(ram_w8_l2048_id0_3_0_wdata),
    .ram_w8_l2048_id0_3_0_wenable(ram_w8_l2048_id0_3_0_wenable),
    .ram_w8_l2048_id0_3_0_enable(ram_w8_l2048_id0_3_0_enable),
    .ram_w8_l2048_id0_3_1_addr(ram_w8_l2048_id0_3_1_addr),
    .ram_w8_l2048_id0_3_1_rdata(ram_w8_l2048_id0_3_1_rdata),
    .ram_w8_l2048_id0_3_1_wdata(ram_w8_l2048_id0_3_1_wdata),
    .ram_w8_l2048_id0_3_1_wenable(ram_w8_l2048_id0_3_1_wenable),
    .ram_w8_l2048_id0_3_1_enable(ram_w8_l2048_id0_3_1_enable)
  );

  wire [9-1:0] ram_w8_l2048_id1_0_0_addr;
  wire [8-1:0] ram_w8_l2048_id1_0_0_rdata;
  wire [8-1:0] ram_w8_l2048_id1_0_0_wdata;
  wire ram_w8_l2048_id1_0_0_wenable;
  wire ram_w8_l2048_id1_0_0_enable;
  wire [9-1:0] ram_w8_l2048_id1_0_1_addr;
  wire [8-1:0] ram_w8_l2048_id1_0_1_rdata;
  wire [8-1:0] ram_w8_l2048_id1_0_1_wdata;
  wire ram_w8_l2048_id1_0_1_wenable;
  wire ram_w8_l2048_id1_0_1_enable;
  assign ram_w8_l2048_id1_0_1_wdata = 'hx;
  assign ram_w8_l2048_id1_0_1_wenable = 0;

  ram_w8_l2048_id1_0
  inst_ram_w8_l2048_id1_0
  (
    .CLK(CLK),
    .ram_w8_l2048_id1_0_0_addr(ram_w8_l2048_id1_0_0_addr),
    .ram_w8_l2048_id1_0_0_rdata(ram_w8_l2048_id1_0_0_rdata),
    .ram_w8_l2048_id1_0_0_wdata(ram_w8_l2048_id1_0_0_wdata),
    .ram_w8_l2048_id1_0_0_wenable(ram_w8_l2048_id1_0_0_wenable),
    .ram_w8_l2048_id1_0_0_enable(ram_w8_l2048_id1_0_0_enable),
    .ram_w8_l2048_id1_0_1_addr(ram_w8_l2048_id1_0_1_addr),
    .ram_w8_l2048_id1_0_1_rdata(ram_w8_l2048_id1_0_1_rdata),
    .ram_w8_l2048_id1_0_1_wdata(ram_w8_l2048_id1_0_1_wdata),
    .ram_w8_l2048_id1_0_1_wenable(ram_w8_l2048_id1_0_1_wenable),
    .ram_w8_l2048_id1_0_1_enable(ram_w8_l2048_id1_0_1_enable)
  );

  wire [9-1:0] ram_w8_l2048_id1_1_0_addr;
  wire [8-1:0] ram_w8_l2048_id1_1_0_rdata;
  wire [8-1:0] ram_w8_l2048_id1_1_0_wdata;
  wire ram_w8_l2048_id1_1_0_wenable;
  wire ram_w8_l2048_id1_1_0_enable;
  wire [9-1:0] ram_w8_l2048_id1_1_1_addr;
  wire [8-1:0] ram_w8_l2048_id1_1_1_rdata;
  wire [8-1:0] ram_w8_l2048_id1_1_1_wdata;
  wire ram_w8_l2048_id1_1_1_wenable;
  wire ram_w8_l2048_id1_1_1_enable;
  assign ram_w8_l2048_id1_1_1_wdata = 'hx;
  assign ram_w8_l2048_id1_1_1_wenable = 0;

  ram_w8_l2048_id1_1
  inst_ram_w8_l2048_id1_1
  (
    .CLK(CLK),
    .ram_w8_l2048_id1_1_0_addr(ram_w8_l2048_id1_1_0_addr),
    .ram_w8_l2048_id1_1_0_rdata(ram_w8_l2048_id1_1_0_rdata),
    .ram_w8_l2048_id1_1_0_wdata(ram_w8_l2048_id1_1_0_wdata),
    .ram_w8_l2048_id1_1_0_wenable(ram_w8_l2048_id1_1_0_wenable),
    .ram_w8_l2048_id1_1_0_enable(ram_w8_l2048_id1_1_0_enable),
    .ram_w8_l2048_id1_1_1_addr(ram_w8_l2048_id1_1_1_addr),
    .ram_w8_l2048_id1_1_1_rdata(ram_w8_l2048_id1_1_1_rdata),
    .ram_w8_l2048_id1_1_1_wdata(ram_w8_l2048_id1_1_1_wdata),
    .ram_w8_l2048_id1_1_1_wenable(ram_w8_l2048_id1_1_1_wenable),
    .ram_w8_l2048_id1_1_1_enable(ram_w8_l2048_id1_1_1_enable)
  );

  wire [9-1:0] ram_w8_l2048_id1_2_0_addr;
  wire [8-1:0] ram_w8_l2048_id1_2_0_rdata;
  wire [8-1:0] ram_w8_l2048_id1_2_0_wdata;
  wire ram_w8_l2048_id1_2_0_wenable;
  wire ram_w8_l2048_id1_2_0_enable;
  wire [9-1:0] ram_w8_l2048_id1_2_1_addr;
  wire [8-1:0] ram_w8_l2048_id1_2_1_rdata;
  wire [8-1:0] ram_w8_l2048_id1_2_1_wdata;
  wire ram_w8_l2048_id1_2_1_wenable;
  wire ram_w8_l2048_id1_2_1_enable;
  assign ram_w8_l2048_id1_2_1_wdata = 'hx;
  assign ram_w8_l2048_id1_2_1_wenable = 0;

  ram_w8_l2048_id1_2
  inst_ram_w8_l2048_id1_2
  (
    .CLK(CLK),
    .ram_w8_l2048_id1_2_0_addr(ram_w8_l2048_id1_2_0_addr),
    .ram_w8_l2048_id1_2_0_rdata(ram_w8_l2048_id1_2_0_rdata),
    .ram_w8_l2048_id1_2_0_wdata(ram_w8_l2048_id1_2_0_wdata),
    .ram_w8_l2048_id1_2_0_wenable(ram_w8_l2048_id1_2_0_wenable),
    .ram_w8_l2048_id1_2_0_enable(ram_w8_l2048_id1_2_0_enable),
    .ram_w8_l2048_id1_2_1_addr(ram_w8_l2048_id1_2_1_addr),
    .ram_w8_l2048_id1_2_1_rdata(ram_w8_l2048_id1_2_1_rdata),
    .ram_w8_l2048_id1_2_1_wdata(ram_w8_l2048_id1_2_1_wdata),
    .ram_w8_l2048_id1_2_1_wenable(ram_w8_l2048_id1_2_1_wenable),
    .ram_w8_l2048_id1_2_1_enable(ram_w8_l2048_id1_2_1_enable)
  );

  wire [9-1:0] ram_w8_l2048_id1_3_0_addr;
  wire [8-1:0] ram_w8_l2048_id1_3_0_rdata;
  wire [8-1:0] ram_w8_l2048_id1_3_0_wdata;
  wire ram_w8_l2048_id1_3_0_wenable;
  wire ram_w8_l2048_id1_3_0_enable;
  wire [9-1:0] ram_w8_l2048_id1_3_1_addr;
  wire [8-1:0] ram_w8_l2048_id1_3_1_rdata;
  wire [8-1:0] ram_w8_l2048_id1_3_1_wdata;
  wire ram_w8_l2048_id1_3_1_wenable;
  wire ram_w8_l2048_id1_3_1_enable;
  assign ram_w8_l2048_id1_3_1_wdata = 'hx;
  assign ram_w8_l2048_id1_3_1_wenable = 0;

  ram_w8_l2048_id1_3
  inst_ram_w8_l2048_id1_3
  (
    .CLK(CLK),
    .ram_w8_l2048_id1_3_0_addr(ram_w8_l2048_id1_3_0_addr),
    .ram_w8_l2048_id1_3_0_rdata(ram_w8_l2048_id1_3_0_rdata),
    .ram_w8_l2048_id1_3_0_wdata(ram_w8_l2048_id1_3_0_wdata),
    .ram_w8_l2048_id1_3_0_wenable(ram_w8_l2048_id1_3_0_wenable),
    .ram_w8_l2048_id1_3_0_enable(ram_w8_l2048_id1_3_0_enable),
    .ram_w8_l2048_id1_3_1_addr(ram_w8_l2048_id1_3_1_addr),
    .ram_w8_l2048_id1_3_1_rdata(ram_w8_l2048_id1_3_1_rdata),
    .ram_w8_l2048_id1_3_1_wdata(ram_w8_l2048_id1_3_1_wdata),
    .ram_w8_l2048_id1_3_1_wenable(ram_w8_l2048_id1_3_1_wenable),
    .ram_w8_l2048_id1_3_1_enable(ram_w8_l2048_id1_3_1_enable)
  );

  wire [8-1:0] cparam_conv2d_24_act_num_col;
  wire [8-1:0] cparam_conv2d_24_act_num_row;
  wire [10-1:0] cparam_conv2d_24_filter_num_och;
  wire [1-1:0] cparam_conv2d_24_bias_scala;
  wire [10-1:0] cparam_conv2d_24_bias_num;
  wire [1-1:0] cparam_conv2d_24_scale_scala;
  wire [1-1:0] cparam_conv2d_24_scale_num;
  wire [1-1:0] cparam_conv2d_24_vshamt_mul_scala;
  wire [1-1:0] cparam_conv2d_24_vshamt_mul_num;
  wire [1-1:0] cparam_conv2d_24_vshamt_sum_scala;
  wire [1-1:0] cparam_conv2d_24_vshamt_sum_num;
  wire [1-1:0] cparam_conv2d_24_vshamt_out_scala;
  wire [1-1:0] cparam_conv2d_24_vshamt_out_num;
  wire [1-1:0] cparam_conv2d_24_cshamt_mul_value;
  wire [1-1:0] cparam_conv2d_24_cshamt_sum_value;
  wire [5-1:0] cparam_conv2d_24_cshamt_out_value;
  wire [1-1:0] cparam_conv2d_24_act_func_index;
  wire [8-1:0] cparam_conv2d_24_out_num_col;
  wire [8-1:0] cparam_conv2d_24_out_num_row;
  wire [1-1:0] cparam_conv2d_24_pad_col_left;
  wire [1-1:0] cparam_conv2d_24_pad_row_top;
  wire [8-1:0] cparam_conv2d_24_max_col_count;
  wire [8-1:0] cparam_conv2d_24_max_row_count;
  wire [1-1:0] cparam_conv2d_24_max_bat_count;
  wire [9-1:0] cparam_conv2d_24_max_och_count;
  wire [5-1:0] cparam_conv2d_24_och_count_step;
  wire [1-1:0] cparam_conv2d_24_dma_flag_conds_0;
  wire [1-1:0] cparam_conv2d_24_dma_flag_conds_1;
  wire [1-1:0] cparam_conv2d_24_dma_flag_conds_2;
  wire signed [32-1:0] cparam_conv2d_24_act_offset_values_0;
  wire signed [32-1:0] cparam_conv2d_24_act_offset_values_1;
  wire signed [32-1:0] cparam_conv2d_24_act_offset_values_2;
  wire [14-1:0] cparam_conv2d_24_act_row_step;
  wire [20-1:0] cparam_conv2d_24_act_bat_step;
  wire [14-1:0] cparam_conv2d_24_act_read_size;
  wire [10-1:0] cparam_conv2d_24_act_read_block;
  wire [13-1:0] cparam_conv2d_24_act_read_step;
  wire [15-1:0] cparam_conv2d_24_filter_base_step;
  wire [15-1:0] cparam_conv2d_24_filter_read_size;
  wire [10-1:0] cparam_conv2d_24_filter_read_block;
  wire [12-1:0] cparam_conv2d_24_filter_read_step;
  wire [1-1:0] cparam_conv2d_24_out_offset_values_0;
  wire [10-1:0] cparam_conv2d_24_out_col_step;
  wire [14-1:0] cparam_conv2d_24_out_row_step;
  wire [22-1:0] cparam_conv2d_24_out_bat_step;
  wire [5-1:0] cparam_conv2d_24_out_och_step;
  wire [5-1:0] cparam_conv2d_24_out_write_size;
  wire [5-1:0] cparam_conv2d_24_out_write_size_res;
  wire [1-1:0] cparam_conv2d_24_out_write_block;
  wire [1-1:0] cparam_conv2d_24_keep_filter;
  wire [1-1:0] cparam_conv2d_24_keep_input;
  wire [1-1:0] cparam_conv2d_24_data_stationary;
  wire [5-1:0] cparam_conv2d_24_stream_num_ops;
  wire [5-1:0] cparam_conv2d_24_stream_num_ops_res;
  wire [5-1:0] cparam_conv2d_24_stream_num_ops_par;
  wire [5-1:0] cparam_conv2d_24_stream_num_ops_res_par;
  wire [10-1:0] cparam_conv2d_24_stream_reduce_size;
  wire [10-1:0] cparam_conv2d_24_stream_aligned_reduce_size;
  wire [1-1:0] cparam_conv2d_24_stream_omit_mask;
  wire [2-1:0] cparam_conv2d_24_col_select_initval;
  wire [1-1:0] cparam_conv2d_24_stride_col_par_col;
  wire [1-1:0] cparam_conv2d_24_stride_row_par_row;
  wire [1-1:0] cparam_conv2d_24_stride_col_mod_filter_num;
  wire [2-1:0] cparam_conv2d_24_filter_num_col_minus_stride_col_mod;
  wire [1-1:0] cparam_conv2d_24_inc_act_laddr_conds_0;
  wire [1-1:0] cparam_conv2d_24_inc_act_laddr_conds_1;
  wire [1-1:0] cparam_conv2d_24_inc_act_laddr_conds_2;
  wire [1-1:0] cparam_conv2d_24_inc_act_laddr_conds_3;
  wire [1-1:0] cparam_conv2d_24_inc_act_laddr_conds_4;
  wire [1-1:0] cparam_conv2d_24_inc_act_laddr_conds_5;
  wire [1-1:0] cparam_conv2d_24_inc_act_laddr_conds_6;
  wire [1-1:0] cparam_conv2d_24_inc_act_laddr_conds_7;
  wire [1-1:0] cparam_conv2d_24_inc_act_laddr_conds_8;
  wire [1-1:0] cparam_conv2d_24_inc_act_laddr_conds_9;
  wire [1-1:0] cparam_conv2d_24_inc_act_laddr_conds_10;
  wire [1-1:0] cparam_conv2d_24_inc_act_laddr_conds_11;
  wire [1-1:0] cparam_conv2d_24_inc_act_laddr_conds_12;
  wire [1-1:0] cparam_conv2d_24_inc_act_laddr_conds_13;
  wire [1-1:0] cparam_conv2d_24_inc_act_laddr_conds_14;
  wire [1-1:0] cparam_conv2d_24_inc_act_laddr_conds_15;
  wire [1-1:0] cparam_conv2d_24_inc_act_laddr_conds_16;
  wire [1-1:0] cparam_conv2d_24_inc_act_laddr_conds_17;
  wire [1-1:0] cparam_conv2d_24_inc_act_laddr_conds_18;
  wire [1-1:0] cparam_conv2d_24_inc_act_laddr_conds_19;
  wire [1-1:0] cparam_conv2d_24_inc_act_laddr_conds_20;
  wire [1-1:0] cparam_conv2d_24_inc_act_laddr_conds_21;
  wire [1-1:0] cparam_conv2d_24_inc_act_laddr_conds_22;
  wire [1-1:0] cparam_conv2d_24_inc_act_laddr_conds_23;
  wire [1-1:0] cparam_conv2d_24_inc_act_laddr_conds_24;
  wire [1-1:0] cparam_conv2d_24_inc_act_laddr_conds_25;
  wire [1-1:0] cparam_conv2d_24_inc_act_laddr_conds_26;
  wire [1-1:0] cparam_conv2d_24_inc_act_laddr_small;
  wire [10-1:0] cparam_conv2d_24_inc_act_laddr_large;
  wire [10-1:0] cparam_conv2d_24_inc_out_laddr_col;
  wire [1-1:0] cparam_conv2d_24_stream_act_local_small_offset;
  wire signed [11-1:0] cparam_conv2d_24_stream_act_local_large_offset;
  wire [1-1:0] cparam_conv2d_24_stream_act_local_small_flags_0;
  wire [1-1:0] cparam_conv2d_24_stream_act_local_small_flags_1;
  wire [1-1:0] cparam_conv2d_24_stream_act_local_small_flags_2;
  wire [1-1:0] cparam_conv2d_24_stream_act_local_large_flags_0;
  wire [1-1:0] cparam_conv2d_24_stream_act_local_large_flags_1;
  wire [1-1:0] cparam_conv2d_24_stream_act_local_large_flags_2;
  wire [1-1:0] cparam_conv2d_24_inc_sync_out;
  wire [1-1:0] cparam_conv2d_24_inc_sync_out_res;
  reg [3-1:0] conv2d_24_control_param_index;
  assign cparam_conv2d_24_act_num_col = (conv2d_24_control_param_index == 0)? 32'he0 : 
                                        (conv2d_24_control_param_index == 1)? 32'h70 : 
                                        (conv2d_24_control_param_index == 2)? 32'h38 : 
                                        (conv2d_24_control_param_index == 3)? 32'h38 : 
                                        (conv2d_24_control_param_index == 4)? 32'h1c : 
                                        (conv2d_24_control_param_index == 5)? 32'h1c : 
                                        (conv2d_24_control_param_index == 6)? 32'he : 32'he;
  assign cparam_conv2d_24_act_num_row = (conv2d_24_control_param_index == 0)? 32'he0 : 
                                        (conv2d_24_control_param_index == 1)? 32'h70 : 
                                        (conv2d_24_control_param_index == 2)? 32'h38 : 
                                        (conv2d_24_control_param_index == 3)? 32'h38 : 
                                        (conv2d_24_control_param_index == 4)? 32'h1c : 
                                        (conv2d_24_control_param_index == 5)? 32'h1c : 
                                        (conv2d_24_control_param_index == 6)? 32'he : 32'he;
  assign cparam_conv2d_24_filter_num_och = (conv2d_24_control_param_index == 0)? 32'h40 : 
                                           (conv2d_24_control_param_index == 1)? 32'h80 : 
                                           (conv2d_24_control_param_index == 2)? 32'h100 : 
                                           (conv2d_24_control_param_index == 3)? 32'h100 : 
                                           (conv2d_24_control_param_index == 4)? 32'h200 : 
                                           (conv2d_24_control_param_index == 5)? 32'h200 : 
                                           (conv2d_24_control_param_index == 6)? 32'h200 : 32'h200;
  assign cparam_conv2d_24_bias_scala = (conv2d_24_control_param_index == 0)? 32'h0 : 
                                       (conv2d_24_control_param_index == 1)? 32'h0 : 
                                       (conv2d_24_control_param_index == 2)? 32'h0 : 
                                       (conv2d_24_control_param_index == 3)? 32'h0 : 
                                       (conv2d_24_control_param_index == 4)? 32'h0 : 
                                       (conv2d_24_control_param_index == 5)? 32'h0 : 
                                       (conv2d_24_control_param_index == 6)? 32'h0 : 32'h0;
  assign cparam_conv2d_24_bias_num = (conv2d_24_control_param_index == 0)? 32'h40 : 
                                     (conv2d_24_control_param_index == 1)? 32'h80 : 
                                     (conv2d_24_control_param_index == 2)? 32'h100 : 
                                     (conv2d_24_control_param_index == 3)? 32'h100 : 
                                     (conv2d_24_control_param_index == 4)? 32'h200 : 
                                     (conv2d_24_control_param_index == 5)? 32'h200 : 
                                     (conv2d_24_control_param_index == 6)? 32'h200 : 32'h200;
  assign cparam_conv2d_24_scale_scala = (conv2d_24_control_param_index == 0)? 32'h1 : 
                                        (conv2d_24_control_param_index == 1)? 32'h1 : 
                                        (conv2d_24_control_param_index == 2)? 32'h1 : 
                                        (conv2d_24_control_param_index == 3)? 32'h1 : 
                                        (conv2d_24_control_param_index == 4)? 32'h1 : 
                                        (conv2d_24_control_param_index == 5)? 32'h1 : 
                                        (conv2d_24_control_param_index == 6)? 32'h1 : 32'h1;
  assign cparam_conv2d_24_scale_num = (conv2d_24_control_param_index == 0)? 32'h1 : 
                                      (conv2d_24_control_param_index == 1)? 32'h1 : 
                                      (conv2d_24_control_param_index == 2)? 32'h1 : 
                                      (conv2d_24_control_param_index == 3)? 32'h1 : 
                                      (conv2d_24_control_param_index == 4)? 32'h1 : 
                                      (conv2d_24_control_param_index == 5)? 32'h1 : 
                                      (conv2d_24_control_param_index == 6)? 32'h1 : 32'h1;
  assign cparam_conv2d_24_vshamt_mul_scala = (conv2d_24_control_param_index == 0)? 32'h0 : 
                                             (conv2d_24_control_param_index == 1)? 32'h0 : 
                                             (conv2d_24_control_param_index == 2)? 32'h0 : 
                                             (conv2d_24_control_param_index == 3)? 32'h0 : 
                                             (conv2d_24_control_param_index == 4)? 32'h0 : 
                                             (conv2d_24_control_param_index == 5)? 32'h0 : 
                                             (conv2d_24_control_param_index == 6)? 32'h0 : 32'h0;
  assign cparam_conv2d_24_vshamt_mul_num = (conv2d_24_control_param_index == 0)? 32'h0 : 
                                           (conv2d_24_control_param_index == 1)? 32'h0 : 
                                           (conv2d_24_control_param_index == 2)? 32'h0 : 
                                           (conv2d_24_control_param_index == 3)? 32'h0 : 
                                           (conv2d_24_control_param_index == 4)? 32'h0 : 
                                           (conv2d_24_control_param_index == 5)? 32'h0 : 
                                           (conv2d_24_control_param_index == 6)? 32'h0 : 32'h0;
  assign cparam_conv2d_24_vshamt_sum_scala = (conv2d_24_control_param_index == 0)? 32'h0 : 
                                             (conv2d_24_control_param_index == 1)? 32'h0 : 
                                             (conv2d_24_control_param_index == 2)? 32'h0 : 
                                             (conv2d_24_control_param_index == 3)? 32'h0 : 
                                             (conv2d_24_control_param_index == 4)? 32'h0 : 
                                             (conv2d_24_control_param_index == 5)? 32'h0 : 
                                             (conv2d_24_control_param_index == 6)? 32'h0 : 32'h0;
  assign cparam_conv2d_24_vshamt_sum_num = (conv2d_24_control_param_index == 0)? 32'h0 : 
                                           (conv2d_24_control_param_index == 1)? 32'h0 : 
                                           (conv2d_24_control_param_index == 2)? 32'h0 : 
                                           (conv2d_24_control_param_index == 3)? 32'h0 : 
                                           (conv2d_24_control_param_index == 4)? 32'h0 : 
                                           (conv2d_24_control_param_index == 5)? 32'h0 : 
                                           (conv2d_24_control_param_index == 6)? 32'h0 : 32'h0;
  assign cparam_conv2d_24_vshamt_out_scala = (conv2d_24_control_param_index == 0)? 32'h0 : 
                                             (conv2d_24_control_param_index == 1)? 32'h0 : 
                                             (conv2d_24_control_param_index == 2)? 32'h0 : 
                                             (conv2d_24_control_param_index == 3)? 32'h0 : 
                                             (conv2d_24_control_param_index == 4)? 32'h0 : 
                                             (conv2d_24_control_param_index == 5)? 32'h0 : 
                                             (conv2d_24_control_param_index == 6)? 32'h0 : 32'h0;
  assign cparam_conv2d_24_vshamt_out_num = (conv2d_24_control_param_index == 0)? 32'h0 : 
                                           (conv2d_24_control_param_index == 1)? 32'h0 : 
                                           (conv2d_24_control_param_index == 2)? 32'h0 : 
                                           (conv2d_24_control_param_index == 3)? 32'h0 : 
                                           (conv2d_24_control_param_index == 4)? 32'h0 : 
                                           (conv2d_24_control_param_index == 5)? 32'h0 : 
                                           (conv2d_24_control_param_index == 6)? 32'h0 : 32'h0;
  assign cparam_conv2d_24_cshamt_mul_value = (conv2d_24_control_param_index == 0)? 32'h0 : 
                                             (conv2d_24_control_param_index == 1)? 32'h0 : 
                                             (conv2d_24_control_param_index == 2)? 32'h0 : 
                                             (conv2d_24_control_param_index == 3)? 32'h0 : 
                                             (conv2d_24_control_param_index == 4)? 32'h0 : 
                                             (conv2d_24_control_param_index == 5)? 32'h0 : 
                                             (conv2d_24_control_param_index == 6)? 32'h0 : 32'h0;
  assign cparam_conv2d_24_cshamt_sum_value = (conv2d_24_control_param_index == 0)? 32'h0 : 
                                             (conv2d_24_control_param_index == 1)? 32'h0 : 
                                             (conv2d_24_control_param_index == 2)? 32'h0 : 
                                             (conv2d_24_control_param_index == 3)? 32'h0 : 
                                             (conv2d_24_control_param_index == 4)? 32'h0 : 
                                             (conv2d_24_control_param_index == 5)? 32'h0 : 
                                             (conv2d_24_control_param_index == 6)? 32'h0 : 32'h0;
  assign cparam_conv2d_24_cshamt_out_value = (conv2d_24_control_param_index == 0)? 32'h10 : 
                                             (conv2d_24_control_param_index == 1)? 32'he : 
                                             (conv2d_24_control_param_index == 2)? 32'hf : 
                                             (conv2d_24_control_param_index == 3)? 32'hf : 
                                             (conv2d_24_control_param_index == 4)? 32'hd : 
                                             (conv2d_24_control_param_index == 5)? 32'he : 
                                             (conv2d_24_control_param_index == 6)? 32'hf : 32'hf;
  assign cparam_conv2d_24_act_func_index = (conv2d_24_control_param_index == 0)? 32'h0 : 
                                           (conv2d_24_control_param_index == 1)? 32'h0 : 
                                           (conv2d_24_control_param_index == 2)? 32'h0 : 
                                           (conv2d_24_control_param_index == 3)? 32'h0 : 
                                           (conv2d_24_control_param_index == 4)? 32'h0 : 
                                           (conv2d_24_control_param_index == 5)? 32'h0 : 
                                           (conv2d_24_control_param_index == 6)? 32'h0 : 32'h0;
  assign cparam_conv2d_24_out_num_col = (conv2d_24_control_param_index == 0)? 32'he0 : 
                                        (conv2d_24_control_param_index == 1)? 32'h70 : 
                                        (conv2d_24_control_param_index == 2)? 32'h38 : 
                                        (conv2d_24_control_param_index == 3)? 32'h38 : 
                                        (conv2d_24_control_param_index == 4)? 32'h1c : 
                                        (conv2d_24_control_param_index == 5)? 32'h1c : 
                                        (conv2d_24_control_param_index == 6)? 32'he : 32'he;
  assign cparam_conv2d_24_out_num_row = (conv2d_24_control_param_index == 0)? 32'he0 : 
                                        (conv2d_24_control_param_index == 1)? 32'h70 : 
                                        (conv2d_24_control_param_index == 2)? 32'h38 : 
                                        (conv2d_24_control_param_index == 3)? 32'h38 : 
                                        (conv2d_24_control_param_index == 4)? 32'h1c : 
                                        (conv2d_24_control_param_index == 5)? 32'h1c : 
                                        (conv2d_24_control_param_index == 6)? 32'he : 32'he;
  assign cparam_conv2d_24_pad_col_left = (conv2d_24_control_param_index == 0)? 32'h1 : 
                                         (conv2d_24_control_param_index == 1)? 32'h1 : 
                                         (conv2d_24_control_param_index == 2)? 32'h1 : 
                                         (conv2d_24_control_param_index == 3)? 32'h1 : 
                                         (conv2d_24_control_param_index == 4)? 32'h1 : 
                                         (conv2d_24_control_param_index == 5)? 32'h1 : 
                                         (conv2d_24_control_param_index == 6)? 32'h1 : 32'h1;
  assign cparam_conv2d_24_pad_row_top = (conv2d_24_control_param_index == 0)? 32'h1 : 
                                        (conv2d_24_control_param_index == 1)? 32'h1 : 
                                        (conv2d_24_control_param_index == 2)? 32'h1 : 
                                        (conv2d_24_control_param_index == 3)? 32'h1 : 
                                        (conv2d_24_control_param_index == 4)? 32'h1 : 
                                        (conv2d_24_control_param_index == 5)? 32'h1 : 
                                        (conv2d_24_control_param_index == 6)? 32'h1 : 32'h1;
  assign cparam_conv2d_24_max_col_count = (conv2d_24_control_param_index == 0)? 32'hdf : 
                                          (conv2d_24_control_param_index == 1)? 32'h6f : 
                                          (conv2d_24_control_param_index == 2)? 32'h37 : 
                                          (conv2d_24_control_param_index == 3)? 32'h37 : 
                                          (conv2d_24_control_param_index == 4)? 32'h1b : 
                                          (conv2d_24_control_param_index == 5)? 32'h1b : 
                                          (conv2d_24_control_param_index == 6)? 32'hd : 32'hd;
  assign cparam_conv2d_24_max_row_count = (conv2d_24_control_param_index == 0)? 32'hdf : 
                                          (conv2d_24_control_param_index == 1)? 32'h6f : 
                                          (conv2d_24_control_param_index == 2)? 32'h37 : 
                                          (conv2d_24_control_param_index == 3)? 32'h37 : 
                                          (conv2d_24_control_param_index == 4)? 32'h1b : 
                                          (conv2d_24_control_param_index == 5)? 32'h1b : 
                                          (conv2d_24_control_param_index == 6)? 32'hd : 32'hd;
  assign cparam_conv2d_24_max_bat_count = (conv2d_24_control_param_index == 0)? 32'h0 : 
                                          (conv2d_24_control_param_index == 1)? 32'h0 : 
                                          (conv2d_24_control_param_index == 2)? 32'h0 : 
                                          (conv2d_24_control_param_index == 3)? 32'h0 : 
                                          (conv2d_24_control_param_index == 4)? 32'h0 : 
                                          (conv2d_24_control_param_index == 5)? 32'h0 : 
                                          (conv2d_24_control_param_index == 6)? 32'h0 : 32'h0;
  assign cparam_conv2d_24_max_och_count = (conv2d_24_control_param_index == 0)? 32'h3c : 
                                          (conv2d_24_control_param_index == 1)? 32'h78 : 
                                          (conv2d_24_control_param_index == 2)? 32'hf0 : 
                                          (conv2d_24_control_param_index == 3)? 32'hf8 : 
                                          (conv2d_24_control_param_index == 4)? 32'h1f8 : 
                                          (conv2d_24_control_param_index == 5)? 32'h1fc : 
                                          (conv2d_24_control_param_index == 6)? 32'h1fc : 32'h1fc;
  assign cparam_conv2d_24_och_count_step = (conv2d_24_control_param_index == 0)? 32'h4 : 
                                           (conv2d_24_control_param_index == 1)? 32'h8 : 
                                           (conv2d_24_control_param_index == 2)? 32'h10 : 
                                           (conv2d_24_control_param_index == 3)? 32'h8 : 
                                           (conv2d_24_control_param_index == 4)? 32'h8 : 
                                           (conv2d_24_control_param_index == 5)? 32'h4 : 
                                           (conv2d_24_control_param_index == 6)? 32'h4 : 32'h4;
  assign cparam_conv2d_24_dma_flag_conds_0 = (conv2d_24_control_param_index == 0)? 32'h1 : 
                                             (conv2d_24_control_param_index == 1)? 32'h1 : 
                                             (conv2d_24_control_param_index == 2)? 32'h1 : 
                                             (conv2d_24_control_param_index == 3)? 32'h1 : 
                                             (conv2d_24_control_param_index == 4)? 32'h1 : 
                                             (conv2d_24_control_param_index == 5)? 32'h1 : 
                                             (conv2d_24_control_param_index == 6)? 32'h1 : 32'h1;
  assign cparam_conv2d_24_dma_flag_conds_1 = (conv2d_24_control_param_index == 0)? 32'h0 : 
                                             (conv2d_24_control_param_index == 1)? 32'h0 : 
                                             (conv2d_24_control_param_index == 2)? 32'h0 : 
                                             (conv2d_24_control_param_index == 3)? 32'h0 : 
                                             (conv2d_24_control_param_index == 4)? 32'h0 : 
                                             (conv2d_24_control_param_index == 5)? 32'h0 : 
                                             (conv2d_24_control_param_index == 6)? 32'h0 : 32'h0;
  assign cparam_conv2d_24_dma_flag_conds_2 = (conv2d_24_control_param_index == 0)? 32'h0 : 
                                             (conv2d_24_control_param_index == 1)? 32'h0 : 
                                             (conv2d_24_control_param_index == 2)? 32'h0 : 
                                             (conv2d_24_control_param_index == 3)? 32'h0 : 
                                             (conv2d_24_control_param_index == 4)? 32'h0 : 
                                             (conv2d_24_control_param_index == 5)? 32'h0 : 
                                             (conv2d_24_control_param_index == 6)? 32'h0 : 32'h0;
  assign cparam_conv2d_24_act_offset_values_0 = (conv2d_24_control_param_index == 0)? -32'sh380 : 
                                                (conv2d_24_control_param_index == 1)? -32'sh1c00 : 
                                                (conv2d_24_control_param_index == 2)? -32'sh1c00 : 
                                                (conv2d_24_control_param_index == 3)? -32'sh3800 : 
                                                (conv2d_24_control_param_index == 4)? -32'sh1c00 : 
                                                (conv2d_24_control_param_index == 5)? -32'sh3800 : 
                                                (conv2d_24_control_param_index == 6)? -32'sh1c00 : -32'sh1c00;
  assign cparam_conv2d_24_act_offset_values_1 = (conv2d_24_control_param_index == 0)? 32'h0 : 
                                                (conv2d_24_control_param_index == 1)? 32'h0 : 
                                                (conv2d_24_control_param_index == 2)? 32'h0 : 
                                                (conv2d_24_control_param_index == 3)? 32'h0 : 
                                                (conv2d_24_control_param_index == 4)? 32'h0 : 
                                                (conv2d_24_control_param_index == 5)? 32'h0 : 
                                                (conv2d_24_control_param_index == 6)? 32'h0 : 32'h0;
  assign cparam_conv2d_24_act_offset_values_2 = (conv2d_24_control_param_index == 0)? 32'h380 : 
                                                (conv2d_24_control_param_index == 1)? 32'h1c00 : 
                                                (conv2d_24_control_param_index == 2)? 32'h1c00 : 
                                                (conv2d_24_control_param_index == 3)? 32'h3800 : 
                                                (conv2d_24_control_param_index == 4)? 32'h1c00 : 
                                                (conv2d_24_control_param_index == 5)? 32'h3800 : 
                                                (conv2d_24_control_param_index == 6)? 32'h1c00 : 32'h1c00;
  assign cparam_conv2d_24_act_row_step = (conv2d_24_control_param_index == 0)? 32'h380 : 
                                         (conv2d_24_control_param_index == 1)? 32'h1c00 : 
                                         (conv2d_24_control_param_index == 2)? 32'h1c00 : 
                                         (conv2d_24_control_param_index == 3)? 32'h3800 : 
                                         (conv2d_24_control_param_index == 4)? 32'h1c00 : 
                                         (conv2d_24_control_param_index == 5)? 32'h3800 : 
                                         (conv2d_24_control_param_index == 6)? 32'h1c00 : 32'h1c00;
  assign cparam_conv2d_24_act_bat_step = (conv2d_24_control_param_index == 0)? 32'h31000 : 
                                         (conv2d_24_control_param_index == 1)? 32'hc4000 : 
                                         (conv2d_24_control_param_index == 2)? 32'h62000 : 
                                         (conv2d_24_control_param_index == 3)? 32'hc4000 : 
                                         (conv2d_24_control_param_index == 4)? 32'h31000 : 
                                         (conv2d_24_control_param_index == 5)? 32'h62000 : 
                                         (conv2d_24_control_param_index == 6)? 32'h18800 : 32'h18800;
  assign cparam_conv2d_24_act_read_size = (conv2d_24_control_param_index == 0)? 32'h380 : 
                                          (conv2d_24_control_param_index == 1)? 32'h1c00 : 
                                          (conv2d_24_control_param_index == 2)? 32'h1c00 : 
                                          (conv2d_24_control_param_index == 3)? 32'h3800 : 
                                          (conv2d_24_control_param_index == 4)? 32'h1c00 : 
                                          (conv2d_24_control_param_index == 5)? 32'h3800 : 
                                          (conv2d_24_control_param_index == 6)? 32'h1c00 : 32'h1c00;
  assign cparam_conv2d_24_act_read_block = (conv2d_24_control_param_index == 0)? 32'h4 : 
                                           (conv2d_24_control_param_index == 1)? 32'h40 : 
                                           (conv2d_24_control_param_index == 2)? 32'h80 : 
                                           (conv2d_24_control_param_index == 3)? 32'h100 : 
                                           (conv2d_24_control_param_index == 4)? 32'h100 : 
                                           (conv2d_24_control_param_index == 5)? 32'h200 : 
                                           (conv2d_24_control_param_index == 6)? 32'h200 : 32'h200;
  assign cparam_conv2d_24_act_read_step = (conv2d_24_control_param_index == 0)? 32'h12c : 
                                          (conv2d_24_control_param_index == 1)? 32'h980 : 
                                          (conv2d_24_control_param_index == 2)? 32'h980 : 
                                          (conv2d_24_control_param_index == 3)? 32'h1300 : 
                                          (conv2d_24_control_param_index == 4)? 32'ha00 : 
                                          (conv2d_24_control_param_index == 5)? 32'h1400 : 
                                          (conv2d_24_control_param_index == 6)? 32'ha00 : 32'ha00;
  assign cparam_conv2d_24_filter_base_step = (conv2d_24_control_param_index == 0)? 32'h90 : 
                                             (conv2d_24_control_param_index == 1)? 32'h1200 : 
                                             (conv2d_24_control_param_index == 2)? 32'h4800 : 
                                             (conv2d_24_control_param_index == 3)? 32'h4800 : 
                                             (conv2d_24_control_param_index == 4)? 32'h4800 : 
                                             (conv2d_24_control_param_index == 5)? 32'h4800 : 
                                             (conv2d_24_control_param_index == 6)? 32'h4800 : 32'h4800;
  assign cparam_conv2d_24_filter_read_size = (conv2d_24_control_param_index == 0)? 32'h90 : 
                                             (conv2d_24_control_param_index == 1)? 32'h1200 : 
                                             (conv2d_24_control_param_index == 2)? 32'h4800 : 
                                             (conv2d_24_control_param_index == 3)? 32'h4800 : 
                                             (conv2d_24_control_param_index == 4)? 32'h4800 : 
                                             (conv2d_24_control_param_index == 5)? 32'h4800 : 
                                             (conv2d_24_control_param_index == 6)? 32'h4800 : 32'h4800;
  assign cparam_conv2d_24_filter_read_block = (conv2d_24_control_param_index == 0)? 32'h4 : 
                                              (conv2d_24_control_param_index == 1)? 32'h40 : 
                                              (conv2d_24_control_param_index == 2)? 32'h80 : 
                                              (conv2d_24_control_param_index == 3)? 32'h100 : 
                                              (conv2d_24_control_param_index == 4)? 32'h100 : 
                                              (conv2d_24_control_param_index == 5)? 32'h200 : 
                                              (conv2d_24_control_param_index == 6)? 32'h200 : 32'h200;
  assign cparam_conv2d_24_filter_read_step = (conv2d_24_control_param_index == 0)? 32'h10 : 
                                             (conv2d_24_control_param_index == 1)? 32'h200 : 
                                             (conv2d_24_control_param_index == 2)? 32'h800 : 
                                             (conv2d_24_control_param_index == 3)? 32'h800 : 
                                             (conv2d_24_control_param_index == 4)? 32'h800 : 
                                             (conv2d_24_control_param_index == 5)? 32'h800 : 
                                             (conv2d_24_control_param_index == 6)? 32'h800 : 32'h800;
  assign cparam_conv2d_24_out_offset_values_0 = (conv2d_24_control_param_index == 0)? 32'h0 : 
                                                (conv2d_24_control_param_index == 1)? 32'h0 : 
                                                (conv2d_24_control_param_index == 2)? 32'h0 : 
                                                (conv2d_24_control_param_index == 3)? 32'h0 : 
                                                (conv2d_24_control_param_index == 4)? 32'h0 : 
                                                (conv2d_24_control_param_index == 5)? 32'h0 : 
                                                (conv2d_24_control_param_index == 6)? 32'h0 : 32'h0;
  assign cparam_conv2d_24_out_col_step = (conv2d_24_control_param_index == 0)? 32'h40 : 
                                         (conv2d_24_control_param_index == 1)? 32'h80 : 
                                         (conv2d_24_control_param_index == 2)? 32'h100 : 
                                         (conv2d_24_control_param_index == 3)? 32'h100 : 
                                         (conv2d_24_control_param_index == 4)? 32'h200 : 
                                         (conv2d_24_control_param_index == 5)? 32'h200 : 
                                         (conv2d_24_control_param_index == 6)? 32'h200 : 32'h200;
  assign cparam_conv2d_24_out_row_step = (conv2d_24_control_param_index == 0)? 32'h3800 : 
                                         (conv2d_24_control_param_index == 1)? 32'h3800 : 
                                         (conv2d_24_control_param_index == 2)? 32'h3800 : 
                                         (conv2d_24_control_param_index == 3)? 32'h3800 : 
                                         (conv2d_24_control_param_index == 4)? 32'h3800 : 
                                         (conv2d_24_control_param_index == 5)? 32'h3800 : 
                                         (conv2d_24_control_param_index == 6)? 32'h1c00 : 32'h1c00;
  assign cparam_conv2d_24_out_bat_step = (conv2d_24_control_param_index == 0)? 32'h310000 : 
                                         (conv2d_24_control_param_index == 1)? 32'h188000 : 
                                         (conv2d_24_control_param_index == 2)? 32'hc4000 : 
                                         (conv2d_24_control_param_index == 3)? 32'hc4000 : 
                                         (conv2d_24_control_param_index == 4)? 32'h62000 : 
                                         (conv2d_24_control_param_index == 5)? 32'h62000 : 
                                         (conv2d_24_control_param_index == 6)? 32'h18800 : 32'h18800;
  assign cparam_conv2d_24_out_och_step = (conv2d_24_control_param_index == 0)? 32'h4 : 
                                         (conv2d_24_control_param_index == 1)? 32'h8 : 
                                         (conv2d_24_control_param_index == 2)? 32'h10 : 
                                         (conv2d_24_control_param_index == 3)? 32'h8 : 
                                         (conv2d_24_control_param_index == 4)? 32'h8 : 
                                         (conv2d_24_control_param_index == 5)? 32'h4 : 
                                         (conv2d_24_control_param_index == 6)? 32'h4 : 32'h4;
  assign cparam_conv2d_24_out_write_size = (conv2d_24_control_param_index == 0)? 32'h4 : 
                                           (conv2d_24_control_param_index == 1)? 32'h8 : 
                                           (conv2d_24_control_param_index == 2)? 32'h10 : 
                                           (conv2d_24_control_param_index == 3)? 32'h8 : 
                                           (conv2d_24_control_param_index == 4)? 32'h8 : 
                                           (conv2d_24_control_param_index == 5)? 32'h4 : 
                                           (conv2d_24_control_param_index == 6)? 32'h4 : 32'h4;
  assign cparam_conv2d_24_out_write_size_res = (conv2d_24_control_param_index == 0)? 32'h4 : 
                                               (conv2d_24_control_param_index == 1)? 32'h8 : 
                                               (conv2d_24_control_param_index == 2)? 32'h10 : 
                                               (conv2d_24_control_param_index == 3)? 32'h8 : 
                                               (conv2d_24_control_param_index == 4)? 32'h8 : 
                                               (conv2d_24_control_param_index == 5)? 32'h4 : 
                                               (conv2d_24_control_param_index == 6)? 32'h4 : 32'h4;
  assign cparam_conv2d_24_out_write_block = (conv2d_24_control_param_index == 0)? 32'h0 : 
                                            (conv2d_24_control_param_index == 1)? 32'h0 : 
                                            (conv2d_24_control_param_index == 2)? 32'h0 : 
                                            (conv2d_24_control_param_index == 3)? 32'h0 : 
                                            (conv2d_24_control_param_index == 4)? 32'h0 : 
                                            (conv2d_24_control_param_index == 5)? 32'h0 : 
                                            (conv2d_24_control_param_index == 6)? 32'h0 : 32'h0;
  assign cparam_conv2d_24_keep_filter = (conv2d_24_control_param_index == 0)? 32'h0 : 
                                        (conv2d_24_control_param_index == 1)? 32'h0 : 
                                        (conv2d_24_control_param_index == 2)? 32'h0 : 
                                        (conv2d_24_control_param_index == 3)? 32'h0 : 
                                        (conv2d_24_control_param_index == 4)? 32'h0 : 
                                        (conv2d_24_control_param_index == 5)? 32'h0 : 
                                        (conv2d_24_control_param_index == 6)? 32'h0 : 32'h0;
  assign cparam_conv2d_24_keep_input = (conv2d_24_control_param_index == 0)? 32'h0 : 
                                       (conv2d_24_control_param_index == 1)? 32'h0 : 
                                       (conv2d_24_control_param_index == 2)? 32'h0 : 
                                       (conv2d_24_control_param_index == 3)? 32'h0 : 
                                       (conv2d_24_control_param_index == 4)? 32'h0 : 
                                       (conv2d_24_control_param_index == 5)? 32'h0 : 
                                       (conv2d_24_control_param_index == 6)? 32'h1 : 32'h1;
  assign cparam_conv2d_24_data_stationary = (conv2d_24_control_param_index == 0)? 32'h0 : 
                                            (conv2d_24_control_param_index == 1)? 32'h0 : 
                                            (conv2d_24_control_param_index == 2)? 32'h0 : 
                                            (conv2d_24_control_param_index == 3)? 32'h0 : 
                                            (conv2d_24_control_param_index == 4)? 32'h0 : 
                                            (conv2d_24_control_param_index == 5)? 32'h0 : 
                                            (conv2d_24_control_param_index == 6)? 32'h0 : 32'h0;
  assign cparam_conv2d_24_stream_num_ops = (conv2d_24_control_param_index == 0)? 32'h4 : 
                                           (conv2d_24_control_param_index == 1)? 32'h8 : 
                                           (conv2d_24_control_param_index == 2)? 32'h10 : 
                                           (conv2d_24_control_param_index == 3)? 32'h8 : 
                                           (conv2d_24_control_param_index == 4)? 32'h8 : 
                                           (conv2d_24_control_param_index == 5)? 32'h4 : 
                                           (conv2d_24_control_param_index == 6)? 32'h4 : 32'h4;
  assign cparam_conv2d_24_stream_num_ops_res = (conv2d_24_control_param_index == 0)? 32'h4 : 
                                               (conv2d_24_control_param_index == 1)? 32'h8 : 
                                               (conv2d_24_control_param_index == 2)? 32'h10 : 
                                               (conv2d_24_control_param_index == 3)? 32'h8 : 
                                               (conv2d_24_control_param_index == 4)? 32'h8 : 
                                               (conv2d_24_control_param_index == 5)? 32'h4 : 
                                               (conv2d_24_control_param_index == 6)? 32'h4 : 32'h4;
  assign cparam_conv2d_24_stream_num_ops_par = (conv2d_24_control_param_index == 0)? 32'h4 : 
                                               (conv2d_24_control_param_index == 1)? 32'h8 : 
                                               (conv2d_24_control_param_index == 2)? 32'h10 : 
                                               (conv2d_24_control_param_index == 3)? 32'h8 : 
                                               (conv2d_24_control_param_index == 4)? 32'h8 : 
                                               (conv2d_24_control_param_index == 5)? 32'h4 : 
                                               (conv2d_24_control_param_index == 6)? 32'h4 : 32'h4;
  assign cparam_conv2d_24_stream_num_ops_res_par = (conv2d_24_control_param_index == 0)? 32'h4 : 
                                                   (conv2d_24_control_param_index == 1)? 32'h8 : 
                                                   (conv2d_24_control_param_index == 2)? 32'h10 : 
                                                   (conv2d_24_control_param_index == 3)? 32'h8 : 
                                                   (conv2d_24_control_param_index == 4)? 32'h8 : 
                                                   (conv2d_24_control_param_index == 5)? 32'h4 : 
                                                   (conv2d_24_control_param_index == 6)? 32'h4 : 32'h4;
  assign cparam_conv2d_24_stream_reduce_size = (conv2d_24_control_param_index == 0)? 32'h3 : 
                                               (conv2d_24_control_param_index == 1)? 32'h40 : 
                                               (conv2d_24_control_param_index == 2)? 32'h80 : 
                                               (conv2d_24_control_param_index == 3)? 32'h100 : 
                                               (conv2d_24_control_param_index == 4)? 32'h100 : 
                                               (conv2d_24_control_param_index == 5)? 32'h200 : 
                                               (conv2d_24_control_param_index == 6)? 32'h200 : 32'h200;
  assign cparam_conv2d_24_stream_aligned_reduce_size = (conv2d_24_control_param_index == 0)? 32'h4 : 
                                                       (conv2d_24_control_param_index == 1)? 32'h40 : 
                                                       (conv2d_24_control_param_index == 2)? 32'h80 : 
                                                       (conv2d_24_control_param_index == 3)? 32'h100 : 
                                                       (conv2d_24_control_param_index == 4)? 32'h100 : 
                                                       (conv2d_24_control_param_index == 5)? 32'h200 : 
                                                       (conv2d_24_control_param_index == 6)? 32'h200 : 32'h200;
  assign cparam_conv2d_24_stream_omit_mask = (conv2d_24_control_param_index == 0)? 32'h0 : 
                                             (conv2d_24_control_param_index == 1)? 32'h0 : 
                                             (conv2d_24_control_param_index == 2)? 32'h0 : 
                                             (conv2d_24_control_param_index == 3)? 32'h0 : 
                                             (conv2d_24_control_param_index == 4)? 32'h0 : 
                                             (conv2d_24_control_param_index == 5)? 32'h0 : 
                                             (conv2d_24_control_param_index == 6)? 32'h0 : 32'h0;
  assign cparam_conv2d_24_col_select_initval = (conv2d_24_control_param_index == 0)? 32'h2 : 
                                               (conv2d_24_control_param_index == 1)? 32'h2 : 
                                               (conv2d_24_control_param_index == 2)? 32'h2 : 
                                               (conv2d_24_control_param_index == 3)? 32'h2 : 
                                               (conv2d_24_control_param_index == 4)? 32'h2 : 
                                               (conv2d_24_control_param_index == 5)? 32'h2 : 
                                               (conv2d_24_control_param_index == 6)? 32'h2 : 32'h2;
  assign cparam_conv2d_24_stride_col_par_col = (conv2d_24_control_param_index == 0)? 32'h1 : 
                                               (conv2d_24_control_param_index == 1)? 32'h1 : 
                                               (conv2d_24_control_param_index == 2)? 32'h1 : 
                                               (conv2d_24_control_param_index == 3)? 32'h1 : 
                                               (conv2d_24_control_param_index == 4)? 32'h1 : 
                                               (conv2d_24_control_param_index == 5)? 32'h1 : 
                                               (conv2d_24_control_param_index == 6)? 32'h1 : 32'h1;
  assign cparam_conv2d_24_stride_row_par_row = (conv2d_24_control_param_index == 0)? 32'h1 : 
                                               (conv2d_24_control_param_index == 1)? 32'h1 : 
                                               (conv2d_24_control_param_index == 2)? 32'h1 : 
                                               (conv2d_24_control_param_index == 3)? 32'h1 : 
                                               (conv2d_24_control_param_index == 4)? 32'h1 : 
                                               (conv2d_24_control_param_index == 5)? 32'h1 : 
                                               (conv2d_24_control_param_index == 6)? 32'h1 : 32'h1;
  assign cparam_conv2d_24_stride_col_mod_filter_num = (conv2d_24_control_param_index == 0)? 32'h1 : 
                                                      (conv2d_24_control_param_index == 1)? 32'h1 : 
                                                      (conv2d_24_control_param_index == 2)? 32'h1 : 
                                                      (conv2d_24_control_param_index == 3)? 32'h1 : 
                                                      (conv2d_24_control_param_index == 4)? 32'h1 : 
                                                      (conv2d_24_control_param_index == 5)? 32'h1 : 
                                                      (conv2d_24_control_param_index == 6)? 32'h1 : 32'h1;
  assign cparam_conv2d_24_filter_num_col_minus_stride_col_mod = (conv2d_24_control_param_index == 0)? 32'h2 : 
                                                                (conv2d_24_control_param_index == 1)? 32'h2 : 
                                                                (conv2d_24_control_param_index == 2)? 32'h2 : 
                                                                (conv2d_24_control_param_index == 3)? 32'h2 : 
                                                                (conv2d_24_control_param_index == 4)? 32'h2 : 
                                                                (conv2d_24_control_param_index == 5)? 32'h2 : 
                                                                (conv2d_24_control_param_index == 6)? 32'h2 : 32'h2;
  assign cparam_conv2d_24_inc_act_laddr_conds_0 = (conv2d_24_control_param_index == 0)? 32'h1 : 
                                                  (conv2d_24_control_param_index == 1)? 32'h1 : 
                                                  (conv2d_24_control_param_index == 2)? 32'h1 : 
                                                  (conv2d_24_control_param_index == 3)? 32'h1 : 
                                                  (conv2d_24_control_param_index == 4)? 32'h1 : 
                                                  (conv2d_24_control_param_index == 5)? 32'h1 : 
                                                  (conv2d_24_control_param_index == 6)? 32'h1 : 32'h1;
  assign cparam_conv2d_24_inc_act_laddr_conds_1 = (conv2d_24_control_param_index == 0)? 32'h0 : 
                                                  (conv2d_24_control_param_index == 1)? 32'h0 : 
                                                  (conv2d_24_control_param_index == 2)? 32'h0 : 
                                                  (conv2d_24_control_param_index == 3)? 32'h0 : 
                                                  (conv2d_24_control_param_index == 4)? 32'h0 : 
                                                  (conv2d_24_control_param_index == 5)? 32'h0 : 
                                                  (conv2d_24_control_param_index == 6)? 32'h0 : 32'h0;
  assign cparam_conv2d_24_inc_act_laddr_conds_2 = (conv2d_24_control_param_index == 0)? 32'h0 : 
                                                  (conv2d_24_control_param_index == 1)? 32'h0 : 
                                                  (conv2d_24_control_param_index == 2)? 32'h0 : 
                                                  (conv2d_24_control_param_index == 3)? 32'h0 : 
                                                  (conv2d_24_control_param_index == 4)? 32'h0 : 
                                                  (conv2d_24_control_param_index == 5)? 32'h0 : 
                                                  (conv2d_24_control_param_index == 6)? 32'h0 : 32'h0;
  assign cparam_conv2d_24_inc_act_laddr_conds_3 = (conv2d_24_control_param_index == 0)? 32'h0 : 
                                                  (conv2d_24_control_param_index == 1)? 32'h0 : 
                                                  (conv2d_24_control_param_index == 2)? 32'h0 : 
                                                  (conv2d_24_control_param_index == 3)? 32'h0 : 
                                                  (conv2d_24_control_param_index == 4)? 32'h0 : 
                                                  (conv2d_24_control_param_index == 5)? 32'h0 : 
                                                  (conv2d_24_control_param_index == 6)? 32'h0 : 32'h0;
  assign cparam_conv2d_24_inc_act_laddr_conds_4 = (conv2d_24_control_param_index == 0)? 32'h1 : 
                                                  (conv2d_24_control_param_index == 1)? 32'h1 : 
                                                  (conv2d_24_control_param_index == 2)? 32'h1 : 
                                                  (conv2d_24_control_param_index == 3)? 32'h1 : 
                                                  (conv2d_24_control_param_index == 4)? 32'h1 : 
                                                  (conv2d_24_control_param_index == 5)? 32'h1 : 
                                                  (conv2d_24_control_param_index == 6)? 32'h1 : 32'h1;
  assign cparam_conv2d_24_inc_act_laddr_conds_5 = (conv2d_24_control_param_index == 0)? 32'h0 : 
                                                  (conv2d_24_control_param_index == 1)? 32'h0 : 
                                                  (conv2d_24_control_param_index == 2)? 32'h0 : 
                                                  (conv2d_24_control_param_index == 3)? 32'h0 : 
                                                  (conv2d_24_control_param_index == 4)? 32'h0 : 
                                                  (conv2d_24_control_param_index == 5)? 32'h0 : 
                                                  (conv2d_24_control_param_index == 6)? 32'h0 : 32'h0;
  assign cparam_conv2d_24_inc_act_laddr_conds_6 = (conv2d_24_control_param_index == 0)? 32'h0 : 
                                                  (conv2d_24_control_param_index == 1)? 32'h0 : 
                                                  (conv2d_24_control_param_index == 2)? 32'h0 : 
                                                  (conv2d_24_control_param_index == 3)? 32'h0 : 
                                                  (conv2d_24_control_param_index == 4)? 32'h0 : 
                                                  (conv2d_24_control_param_index == 5)? 32'h0 : 
                                                  (conv2d_24_control_param_index == 6)? 32'h0 : 32'h0;
  assign cparam_conv2d_24_inc_act_laddr_conds_7 = (conv2d_24_control_param_index == 0)? 32'h0 : 
                                                  (conv2d_24_control_param_index == 1)? 32'h0 : 
                                                  (conv2d_24_control_param_index == 2)? 32'h0 : 
                                                  (conv2d_24_control_param_index == 3)? 32'h0 : 
                                                  (conv2d_24_control_param_index == 4)? 32'h0 : 
                                                  (conv2d_24_control_param_index == 5)? 32'h0 : 
                                                  (conv2d_24_control_param_index == 6)? 32'h0 : 32'h0;
  assign cparam_conv2d_24_inc_act_laddr_conds_8 = (conv2d_24_control_param_index == 0)? 32'h1 : 
                                                  (conv2d_24_control_param_index == 1)? 32'h1 : 
                                                  (conv2d_24_control_param_index == 2)? 32'h1 : 
                                                  (conv2d_24_control_param_index == 3)? 32'h1 : 
                                                  (conv2d_24_control_param_index == 4)? 32'h1 : 
                                                  (conv2d_24_control_param_index == 5)? 32'h1 : 
                                                  (conv2d_24_control_param_index == 6)? 32'h1 : 32'h1;
  assign cparam_conv2d_24_inc_act_laddr_conds_9 = (conv2d_24_control_param_index == 0)? 32'h1 : 
                                                  (conv2d_24_control_param_index == 1)? 32'h1 : 
                                                  (conv2d_24_control_param_index == 2)? 32'h1 : 
                                                  (conv2d_24_control_param_index == 3)? 32'h1 : 
                                                  (conv2d_24_control_param_index == 4)? 32'h1 : 
                                                  (conv2d_24_control_param_index == 5)? 32'h1 : 
                                                  (conv2d_24_control_param_index == 6)? 32'h1 : 32'h1;
  assign cparam_conv2d_24_inc_act_laddr_conds_10 = (conv2d_24_control_param_index == 0)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 1)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 2)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 3)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 4)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 5)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 6)? 32'h0 : 32'h0;
  assign cparam_conv2d_24_inc_act_laddr_conds_11 = (conv2d_24_control_param_index == 0)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 1)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 2)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 3)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 4)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 5)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 6)? 32'h0 : 32'h0;
  assign cparam_conv2d_24_inc_act_laddr_conds_12 = (conv2d_24_control_param_index == 0)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 1)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 2)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 3)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 4)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 5)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 6)? 32'h0 : 32'h0;
  assign cparam_conv2d_24_inc_act_laddr_conds_13 = (conv2d_24_control_param_index == 0)? 32'h1 : 
                                                   (conv2d_24_control_param_index == 1)? 32'h1 : 
                                                   (conv2d_24_control_param_index == 2)? 32'h1 : 
                                                   (conv2d_24_control_param_index == 3)? 32'h1 : 
                                                   (conv2d_24_control_param_index == 4)? 32'h1 : 
                                                   (conv2d_24_control_param_index == 5)? 32'h1 : 
                                                   (conv2d_24_control_param_index == 6)? 32'h1 : 32'h1;
  assign cparam_conv2d_24_inc_act_laddr_conds_14 = (conv2d_24_control_param_index == 0)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 1)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 2)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 3)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 4)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 5)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 6)? 32'h0 : 32'h0;
  assign cparam_conv2d_24_inc_act_laddr_conds_15 = (conv2d_24_control_param_index == 0)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 1)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 2)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 3)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 4)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 5)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 6)? 32'h0 : 32'h0;
  assign cparam_conv2d_24_inc_act_laddr_conds_16 = (conv2d_24_control_param_index == 0)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 1)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 2)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 3)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 4)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 5)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 6)? 32'h0 : 32'h0;
  assign cparam_conv2d_24_inc_act_laddr_conds_17 = (conv2d_24_control_param_index == 0)? 32'h1 : 
                                                   (conv2d_24_control_param_index == 1)? 32'h1 : 
                                                   (conv2d_24_control_param_index == 2)? 32'h1 : 
                                                   (conv2d_24_control_param_index == 3)? 32'h1 : 
                                                   (conv2d_24_control_param_index == 4)? 32'h1 : 
                                                   (conv2d_24_control_param_index == 5)? 32'h1 : 
                                                   (conv2d_24_control_param_index == 6)? 32'h1 : 32'h1;
  assign cparam_conv2d_24_inc_act_laddr_conds_18 = (conv2d_24_control_param_index == 0)? 32'h1 : 
                                                   (conv2d_24_control_param_index == 1)? 32'h1 : 
                                                   (conv2d_24_control_param_index == 2)? 32'h1 : 
                                                   (conv2d_24_control_param_index == 3)? 32'h1 : 
                                                   (conv2d_24_control_param_index == 4)? 32'h1 : 
                                                   (conv2d_24_control_param_index == 5)? 32'h1 : 
                                                   (conv2d_24_control_param_index == 6)? 32'h1 : 32'h1;
  assign cparam_conv2d_24_inc_act_laddr_conds_19 = (conv2d_24_control_param_index == 0)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 1)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 2)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 3)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 4)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 5)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 6)? 32'h0 : 32'h0;
  assign cparam_conv2d_24_inc_act_laddr_conds_20 = (conv2d_24_control_param_index == 0)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 1)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 2)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 3)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 4)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 5)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 6)? 32'h0 : 32'h0;
  assign cparam_conv2d_24_inc_act_laddr_conds_21 = (conv2d_24_control_param_index == 0)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 1)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 2)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 3)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 4)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 5)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 6)? 32'h0 : 32'h0;
  assign cparam_conv2d_24_inc_act_laddr_conds_22 = (conv2d_24_control_param_index == 0)? 32'h1 : 
                                                   (conv2d_24_control_param_index == 1)? 32'h1 : 
                                                   (conv2d_24_control_param_index == 2)? 32'h1 : 
                                                   (conv2d_24_control_param_index == 3)? 32'h1 : 
                                                   (conv2d_24_control_param_index == 4)? 32'h1 : 
                                                   (conv2d_24_control_param_index == 5)? 32'h1 : 
                                                   (conv2d_24_control_param_index == 6)? 32'h1 : 32'h1;
  assign cparam_conv2d_24_inc_act_laddr_conds_23 = (conv2d_24_control_param_index == 0)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 1)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 2)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 3)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 4)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 5)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 6)? 32'h0 : 32'h0;
  assign cparam_conv2d_24_inc_act_laddr_conds_24 = (conv2d_24_control_param_index == 0)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 1)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 2)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 3)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 4)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 5)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 6)? 32'h0 : 32'h0;
  assign cparam_conv2d_24_inc_act_laddr_conds_25 = (conv2d_24_control_param_index == 0)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 1)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 2)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 3)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 4)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 5)? 32'h0 : 
                                                   (conv2d_24_control_param_index == 6)? 32'h0 : 32'h0;
  assign cparam_conv2d_24_inc_act_laddr_conds_26 = (conv2d_24_control_param_index == 0)? 32'h1 : 
                                                   (conv2d_24_control_param_index == 1)? 32'h1 : 
                                                   (conv2d_24_control_param_index == 2)? 32'h1 : 
                                                   (conv2d_24_control_param_index == 3)? 32'h1 : 
                                                   (conv2d_24_control_param_index == 4)? 32'h1 : 
                                                   (conv2d_24_control_param_index == 5)? 32'h1 : 
                                                   (conv2d_24_control_param_index == 6)? 32'h1 : 32'h1;
  assign cparam_conv2d_24_inc_act_laddr_small = (conv2d_24_control_param_index == 0)? 32'h0 : 
                                                (conv2d_24_control_param_index == 1)? 32'h0 : 
                                                (conv2d_24_control_param_index == 2)? 32'h0 : 
                                                (conv2d_24_control_param_index == 3)? 32'h0 : 
                                                (conv2d_24_control_param_index == 4)? 32'h0 : 
                                                (conv2d_24_control_param_index == 5)? 32'h0 : 
                                                (conv2d_24_control_param_index == 6)? 32'h0 : 32'h0;
  assign cparam_conv2d_24_inc_act_laddr_large = (conv2d_24_control_param_index == 0)? 32'h4 : 
                                                (conv2d_24_control_param_index == 1)? 32'h40 : 
                                                (conv2d_24_control_param_index == 2)? 32'h80 : 
                                                (conv2d_24_control_param_index == 3)? 32'h100 : 
                                                (conv2d_24_control_param_index == 4)? 32'h100 : 
                                                (conv2d_24_control_param_index == 5)? 32'h200 : 
                                                (conv2d_24_control_param_index == 6)? 32'h200 : 32'h200;
  assign cparam_conv2d_24_inc_out_laddr_col = (conv2d_24_control_param_index == 0)? 32'h40 : 
                                              (conv2d_24_control_param_index == 1)? 32'h80 : 
                                              (conv2d_24_control_param_index == 2)? 32'h100 : 
                                              (conv2d_24_control_param_index == 3)? 32'h100 : 
                                              (conv2d_24_control_param_index == 4)? 32'h200 : 
                                              (conv2d_24_control_param_index == 5)? 32'h200 : 
                                              (conv2d_24_control_param_index == 6)? 32'h200 : 32'h200;
  assign cparam_conv2d_24_stream_act_local_small_offset = (conv2d_24_control_param_index == 0)? 32'h0 : 
                                                          (conv2d_24_control_param_index == 1)? 32'h0 : 
                                                          (conv2d_24_control_param_index == 2)? 32'h0 : 
                                                          (conv2d_24_control_param_index == 3)? 32'h0 : 
                                                          (conv2d_24_control_param_index == 4)? 32'h0 : 
                                                          (conv2d_24_control_param_index == 5)? 32'h0 : 
                                                          (conv2d_24_control_param_index == 6)? 32'h0 : 32'h0;
  assign cparam_conv2d_24_stream_act_local_large_offset = (conv2d_24_control_param_index == 0)? -32'sh4 : 
                                                          (conv2d_24_control_param_index == 1)? -32'sh40 : 
                                                          (conv2d_24_control_param_index == 2)? -32'sh80 : 
                                                          (conv2d_24_control_param_index == 3)? -32'sh100 : 
                                                          (conv2d_24_control_param_index == 4)? -32'sh100 : 
                                                          (conv2d_24_control_param_index == 5)? -32'sh200 : 
                                                          (conv2d_24_control_param_index == 6)? -32'sh200 : -32'sh200;
  assign cparam_conv2d_24_stream_act_local_small_flags_0 = (conv2d_24_control_param_index == 0)? 32'h0 : 
                                                           (conv2d_24_control_param_index == 1)? 32'h0 : 
                                                           (conv2d_24_control_param_index == 2)? 32'h0 : 
                                                           (conv2d_24_control_param_index == 3)? 32'h0 : 
                                                           (conv2d_24_control_param_index == 4)? 32'h0 : 
                                                           (conv2d_24_control_param_index == 5)? 32'h0 : 
                                                           (conv2d_24_control_param_index == 6)? 32'h0 : 32'h0;
  assign cparam_conv2d_24_stream_act_local_small_flags_1 = (conv2d_24_control_param_index == 0)? 32'h0 : 
                                                           (conv2d_24_control_param_index == 1)? 32'h0 : 
                                                           (conv2d_24_control_param_index == 2)? 32'h0 : 
                                                           (conv2d_24_control_param_index == 3)? 32'h0 : 
                                                           (conv2d_24_control_param_index == 4)? 32'h0 : 
                                                           (conv2d_24_control_param_index == 5)? 32'h0 : 
                                                           (conv2d_24_control_param_index == 6)? 32'h0 : 32'h0;
  assign cparam_conv2d_24_stream_act_local_small_flags_2 = (conv2d_24_control_param_index == 0)? 32'h1 : 
                                                           (conv2d_24_control_param_index == 1)? 32'h1 : 
                                                           (conv2d_24_control_param_index == 2)? 32'h1 : 
                                                           (conv2d_24_control_param_index == 3)? 32'h1 : 
                                                           (conv2d_24_control_param_index == 4)? 32'h1 : 
                                                           (conv2d_24_control_param_index == 5)? 32'h1 : 
                                                           (conv2d_24_control_param_index == 6)? 32'h1 : 32'h1;
  assign cparam_conv2d_24_stream_act_local_large_flags_0 = (conv2d_24_control_param_index == 0)? 32'h0 : 
                                                           (conv2d_24_control_param_index == 1)? 32'h0 : 
                                                           (conv2d_24_control_param_index == 2)? 32'h0 : 
                                                           (conv2d_24_control_param_index == 3)? 32'h0 : 
                                                           (conv2d_24_control_param_index == 4)? 32'h0 : 
                                                           (conv2d_24_control_param_index == 5)? 32'h0 : 
                                                           (conv2d_24_control_param_index == 6)? 32'h0 : 32'h0;
  assign cparam_conv2d_24_stream_act_local_large_flags_1 = (conv2d_24_control_param_index == 0)? 32'h0 : 
                                                           (conv2d_24_control_param_index == 1)? 32'h0 : 
                                                           (conv2d_24_control_param_index == 2)? 32'h0 : 
                                                           (conv2d_24_control_param_index == 3)? 32'h0 : 
                                                           (conv2d_24_control_param_index == 4)? 32'h0 : 
                                                           (conv2d_24_control_param_index == 5)? 32'h0 : 
                                                           (conv2d_24_control_param_index == 6)? 32'h0 : 32'h0;
  assign cparam_conv2d_24_stream_act_local_large_flags_2 = (conv2d_24_control_param_index == 0)? 32'h1 : 
                                                           (conv2d_24_control_param_index == 1)? 32'h1 : 
                                                           (conv2d_24_control_param_index == 2)? 32'h1 : 
                                                           (conv2d_24_control_param_index == 3)? 32'h1 : 
                                                           (conv2d_24_control_param_index == 4)? 32'h1 : 
                                                           (conv2d_24_control_param_index == 5)? 32'h1 : 
                                                           (conv2d_24_control_param_index == 6)? 32'h1 : 32'h1;
  assign cparam_conv2d_24_inc_sync_out = (conv2d_24_control_param_index == 0)? 32'h1 : 
                                         (conv2d_24_control_param_index == 1)? 32'h1 : 
                                         (conv2d_24_control_param_index == 2)? 32'h1 : 
                                         (conv2d_24_control_param_index == 3)? 32'h1 : 
                                         (conv2d_24_control_param_index == 4)? 32'h1 : 
                                         (conv2d_24_control_param_index == 5)? 32'h1 : 
                                         (conv2d_24_control_param_index == 6)? 32'h1 : 32'h1;
  assign cparam_conv2d_24_inc_sync_out_res = (conv2d_24_control_param_index == 0)? 32'h0 : 
                                             (conv2d_24_control_param_index == 1)? 32'h0 : 
                                             (conv2d_24_control_param_index == 2)? 32'h0 : 
                                             (conv2d_24_control_param_index == 3)? 32'h0 : 
                                             (conv2d_24_control_param_index == 4)? 32'h0 : 
                                             (conv2d_24_control_param_index == 5)? 32'h0 : 
                                             (conv2d_24_control_param_index == 6)? 32'h0 : 32'h0;
  wire [8-1:0] cparam_max_pool_serial_26_act_num_col;
  wire [8-1:0] cparam_max_pool_serial_26_act_num_row;
  wire [2-1:0] cparam_max_pool_serial_26_stride_col;
  wire [2-1:0] cparam_max_pool_serial_26_stride_row;
  wire [7-1:0] cparam_max_pool_serial_26_out_num_col;
  wire [7-1:0] cparam_max_pool_serial_26_out_num_row;
  wire [1-1:0] cparam_max_pool_serial_26_pad_col_left;
  wire [1-1:0] cparam_max_pool_serial_26_pad_row_top;
  wire [8-1:0] cparam_max_pool_serial_26_max_col_count;
  wire [8-1:0] cparam_max_pool_serial_26_max_row_count;
  wire [1-1:0] cparam_max_pool_serial_26_max_bat_count;
  wire signed [32-1:0] cparam_max_pool_serial_26_act_offset_values_0;
  wire signed [32-1:0] cparam_max_pool_serial_26_act_offset_values_1;
  wire [15-1:0] cparam_max_pool_serial_26_act_row_step;
  wire [22-1:0] cparam_max_pool_serial_26_act_bat_step;
  wire [14-1:0] cparam_max_pool_serial_26_act_read_size;
  wire [10-1:0] cparam_max_pool_serial_26_act_read_block;
  wire [13-1:0] cparam_max_pool_serial_26_out_row_step;
  wire [20-1:0] cparam_max_pool_serial_26_out_bat_step;
  wire [13-1:0] cparam_max_pool_serial_26_out_write_size;
  wire [10-1:0] cparam_max_pool_serial_26_stream_size;
  wire [1-1:0] cparam_max_pool_serial_26_col_select_initval;
  wire [1-1:0] cparam_max_pool_serial_26_stride_col_mod_ksize;
  wire [2-1:0] cparam_max_pool_serial_26_ksize_col_minus_stride_col_mod;
  wire [1-1:0] cparam_max_pool_serial_26_local_pad_offset;
  wire [11-1:0] cparam_max_pool_serial_26_inc_act_laddr;
  wire [10-1:0] cparam_max_pool_serial_26_inc_out_laddr;
  reg [3-1:0] max_pool_serial_26_control_param_index;
  assign cparam_max_pool_serial_26_act_num_col = (max_pool_serial_26_control_param_index == 0)? 32'he0 : 
                                                 (max_pool_serial_26_control_param_index == 1)? 32'h70 : 
                                                 (max_pool_serial_26_control_param_index == 2)? 32'h38 : 
                                                 (max_pool_serial_26_control_param_index == 3)? 32'h1c : 32'he;
  assign cparam_max_pool_serial_26_act_num_row = (max_pool_serial_26_control_param_index == 0)? 32'he0 : 
                                                 (max_pool_serial_26_control_param_index == 1)? 32'h70 : 
                                                 (max_pool_serial_26_control_param_index == 2)? 32'h38 : 
                                                 (max_pool_serial_26_control_param_index == 3)? 32'h1c : 32'he;
  assign cparam_max_pool_serial_26_stride_col = (max_pool_serial_26_control_param_index == 0)? 32'h2 : 
                                                (max_pool_serial_26_control_param_index == 1)? 32'h2 : 
                                                (max_pool_serial_26_control_param_index == 2)? 32'h2 : 
                                                (max_pool_serial_26_control_param_index == 3)? 32'h2 : 32'h2;
  assign cparam_max_pool_serial_26_stride_row = (max_pool_serial_26_control_param_index == 0)? 32'h2 : 
                                                (max_pool_serial_26_control_param_index == 1)? 32'h2 : 
                                                (max_pool_serial_26_control_param_index == 2)? 32'h2 : 
                                                (max_pool_serial_26_control_param_index == 3)? 32'h2 : 32'h2;
  assign cparam_max_pool_serial_26_out_num_col = (max_pool_serial_26_control_param_index == 0)? 32'h70 : 
                                                 (max_pool_serial_26_control_param_index == 1)? 32'h38 : 
                                                 (max_pool_serial_26_control_param_index == 2)? 32'h1c : 
                                                 (max_pool_serial_26_control_param_index == 3)? 32'he : 32'h7;
  assign cparam_max_pool_serial_26_out_num_row = (max_pool_serial_26_control_param_index == 0)? 32'h70 : 
                                                 (max_pool_serial_26_control_param_index == 1)? 32'h38 : 
                                                 (max_pool_serial_26_control_param_index == 2)? 32'h1c : 
                                                 (max_pool_serial_26_control_param_index == 3)? 32'he : 32'h7;
  assign cparam_max_pool_serial_26_pad_col_left = (max_pool_serial_26_control_param_index == 0)? 32'h0 : 
                                                  (max_pool_serial_26_control_param_index == 1)? 32'h0 : 
                                                  (max_pool_serial_26_control_param_index == 2)? 32'h0 : 
                                                  (max_pool_serial_26_control_param_index == 3)? 32'h0 : 32'h0;
  assign cparam_max_pool_serial_26_pad_row_top = (max_pool_serial_26_control_param_index == 0)? 32'h0 : 
                                                 (max_pool_serial_26_control_param_index == 1)? 32'h0 : 
                                                 (max_pool_serial_26_control_param_index == 2)? 32'h0 : 
                                                 (max_pool_serial_26_control_param_index == 3)? 32'h0 : 32'h0;
  assign cparam_max_pool_serial_26_max_col_count = (max_pool_serial_26_control_param_index == 0)? 32'hdd : 
                                                   (max_pool_serial_26_control_param_index == 1)? 32'h6d : 
                                                   (max_pool_serial_26_control_param_index == 2)? 32'h35 : 
                                                   (max_pool_serial_26_control_param_index == 3)? 32'h19 : 32'hb;
  assign cparam_max_pool_serial_26_max_row_count = (max_pool_serial_26_control_param_index == 0)? 32'hdd : 
                                                   (max_pool_serial_26_control_param_index == 1)? 32'h6d : 
                                                   (max_pool_serial_26_control_param_index == 2)? 32'h35 : 
                                                   (max_pool_serial_26_control_param_index == 3)? 32'h19 : 32'hb;
  assign cparam_max_pool_serial_26_max_bat_count = (max_pool_serial_26_control_param_index == 0)? 32'h0 : 
                                                   (max_pool_serial_26_control_param_index == 1)? 32'h0 : 
                                                   (max_pool_serial_26_control_param_index == 2)? 32'h0 : 
                                                   (max_pool_serial_26_control_param_index == 3)? 32'h0 : 32'h0;
  assign cparam_max_pool_serial_26_act_offset_values_0 = (max_pool_serial_26_control_param_index == 0)? 32'h0 : 
                                                         (max_pool_serial_26_control_param_index == 1)? 32'h0 : 
                                                         (max_pool_serial_26_control_param_index == 2)? 32'h0 : 
                                                         (max_pool_serial_26_control_param_index == 3)? 32'h0 : 32'h0;
  assign cparam_max_pool_serial_26_act_offset_values_1 = (max_pool_serial_26_control_param_index == 0)? 32'h3800 : 
                                                         (max_pool_serial_26_control_param_index == 1)? 32'h3800 : 
                                                         (max_pool_serial_26_control_param_index == 2)? 32'h3800 : 
                                                         (max_pool_serial_26_control_param_index == 3)? 32'h3800 : 32'h1c00;
  assign cparam_max_pool_serial_26_act_row_step = (max_pool_serial_26_control_param_index == 0)? 32'h7000 : 
                                                  (max_pool_serial_26_control_param_index == 1)? 32'h7000 : 
                                                  (max_pool_serial_26_control_param_index == 2)? 32'h7000 : 
                                                  (max_pool_serial_26_control_param_index == 3)? 32'h7000 : 32'h3800;
  assign cparam_max_pool_serial_26_act_bat_step = (max_pool_serial_26_control_param_index == 0)? 32'h310000 : 
                                                  (max_pool_serial_26_control_param_index == 1)? 32'h188000 : 
                                                  (max_pool_serial_26_control_param_index == 2)? 32'hc4000 : 
                                                  (max_pool_serial_26_control_param_index == 3)? 32'h62000 : 32'h18800;
  assign cparam_max_pool_serial_26_act_read_size = (max_pool_serial_26_control_param_index == 0)? 32'h3800 : 
                                                   (max_pool_serial_26_control_param_index == 1)? 32'h3800 : 
                                                   (max_pool_serial_26_control_param_index == 2)? 32'h3800 : 
                                                   (max_pool_serial_26_control_param_index == 3)? 32'h3800 : 32'h1c00;
  assign cparam_max_pool_serial_26_act_read_block = (max_pool_serial_26_control_param_index == 0)? 32'h40 : 
                                                    (max_pool_serial_26_control_param_index == 1)? 32'h80 : 
                                                    (max_pool_serial_26_control_param_index == 2)? 32'h100 : 
                                                    (max_pool_serial_26_control_param_index == 3)? 32'h200 : 32'h200;
  assign cparam_max_pool_serial_26_out_row_step = (max_pool_serial_26_control_param_index == 0)? 32'h1c00 : 
                                                  (max_pool_serial_26_control_param_index == 1)? 32'h1c00 : 
                                                  (max_pool_serial_26_control_param_index == 2)? 32'h1c00 : 
                                                  (max_pool_serial_26_control_param_index == 3)? 32'h1c00 : 32'he00;
  assign cparam_max_pool_serial_26_out_bat_step = (max_pool_serial_26_control_param_index == 0)? 32'hc4000 : 
                                                  (max_pool_serial_26_control_param_index == 1)? 32'h62000 : 
                                                  (max_pool_serial_26_control_param_index == 2)? 32'h31000 : 
                                                  (max_pool_serial_26_control_param_index == 3)? 32'h18800 : 32'h6200;
  assign cparam_max_pool_serial_26_out_write_size = (max_pool_serial_26_control_param_index == 0)? 32'h1c00 : 
                                                    (max_pool_serial_26_control_param_index == 1)? 32'h1c00 : 
                                                    (max_pool_serial_26_control_param_index == 2)? 32'h1c00 : 
                                                    (max_pool_serial_26_control_param_index == 3)? 32'h1c00 : 32'he00;
  assign cparam_max_pool_serial_26_stream_size = (max_pool_serial_26_control_param_index == 0)? 32'h40 : 
                                                 (max_pool_serial_26_control_param_index == 1)? 32'h80 : 
                                                 (max_pool_serial_26_control_param_index == 2)? 32'h100 : 
                                                 (max_pool_serial_26_control_param_index == 3)? 32'h200 : 32'h200;
  assign cparam_max_pool_serial_26_col_select_initval = (max_pool_serial_26_control_param_index == 0)? 32'h0 : 
                                                        (max_pool_serial_26_control_param_index == 1)? 32'h0 : 
                                                        (max_pool_serial_26_control_param_index == 2)? 32'h0 : 
                                                        (max_pool_serial_26_control_param_index == 3)? 32'h0 : 32'h0;
  assign cparam_max_pool_serial_26_stride_col_mod_ksize = (max_pool_serial_26_control_param_index == 0)? 32'h0 : 
                                                          (max_pool_serial_26_control_param_index == 1)? 32'h0 : 
                                                          (max_pool_serial_26_control_param_index == 2)? 32'h0 : 
                                                          (max_pool_serial_26_control_param_index == 3)? 32'h0 : 32'h0;
  assign cparam_max_pool_serial_26_ksize_col_minus_stride_col_mod = (max_pool_serial_26_control_param_index == 0)? 32'h2 : 
                                                                    (max_pool_serial_26_control_param_index == 1)? 32'h2 : 
                                                                    (max_pool_serial_26_control_param_index == 2)? 32'h2 : 
                                                                    (max_pool_serial_26_control_param_index == 3)? 32'h2 : 32'h2;
  assign cparam_max_pool_serial_26_local_pad_offset = (max_pool_serial_26_control_param_index == 0)? 32'h0 : 
                                                      (max_pool_serial_26_control_param_index == 1)? 32'h0 : 
                                                      (max_pool_serial_26_control_param_index == 2)? 32'h0 : 
                                                      (max_pool_serial_26_control_param_index == 3)? 32'h0 : 32'h0;
  assign cparam_max_pool_serial_26_inc_act_laddr = (max_pool_serial_26_control_param_index == 0)? 32'h80 : 
                                                   (max_pool_serial_26_control_param_index == 1)? 32'h100 : 
                                                   (max_pool_serial_26_control_param_index == 2)? 32'h200 : 
                                                   (max_pool_serial_26_control_param_index == 3)? 32'h400 : 32'h400;
  assign cparam_max_pool_serial_26_inc_out_laddr = (max_pool_serial_26_control_param_index == 0)? 32'h40 : 
                                                   (max_pool_serial_26_control_param_index == 1)? 32'h80 : 
                                                   (max_pool_serial_26_control_param_index == 2)? 32'h100 : 
                                                   (max_pool_serial_26_control_param_index == 3)? 32'h200 : 32'h200;
  wire [3-1:0] cparam_avg_pool_serial_52_act_num_col;
  wire [3-1:0] cparam_avg_pool_serial_52_act_num_row;
  wire [1-1:0] cparam_avg_pool_serial_52_stride_col;
  wire [1-1:0] cparam_avg_pool_serial_52_stride_row;
  wire [3-1:0] cparam_avg_pool_serial_52_out_num_col;
  wire [3-1:0] cparam_avg_pool_serial_52_out_num_row;
  wire [1-1:0] cparam_avg_pool_serial_52_pad_col_left;
  wire [1-1:0] cparam_avg_pool_serial_52_pad_row_top;
  wire [3-1:0] cparam_avg_pool_serial_52_max_col_count;
  wire [3-1:0] cparam_avg_pool_serial_52_max_row_count;
  wire [1-1:0] cparam_avg_pool_serial_52_max_bat_count;
  wire signed [32-1:0] cparam_avg_pool_serial_52_act_offset_values_0;
  wire [12-1:0] cparam_avg_pool_serial_52_act_row_step;
  wire [15-1:0] cparam_avg_pool_serial_52_act_bat_step;
  wire [12-1:0] cparam_avg_pool_serial_52_act_read_size;
  wire [10-1:0] cparam_avg_pool_serial_52_act_read_block;
  wire [12-1:0] cparam_avg_pool_serial_52_out_row_step;
  wire [15-1:0] cparam_avg_pool_serial_52_out_bat_step;
  wire [12-1:0] cparam_avg_pool_serial_52_out_write_size;
  wire [10-1:0] cparam_avg_pool_serial_52_stream_size;
  wire [1-1:0] cparam_avg_pool_serial_52_col_select_initval;
  wire [1-1:0] cparam_avg_pool_serial_52_stride_col_mod_ksize;
  wire [1-1:0] cparam_avg_pool_serial_52_ksize_col_minus_stride_col_mod;
  wire [1-1:0] cparam_avg_pool_serial_52_local_pad_offset;
  wire [10-1:0] cparam_avg_pool_serial_52_inc_act_laddr;
  wire [10-1:0] cparam_avg_pool_serial_52_inc_out_laddr;
  assign cparam_avg_pool_serial_52_act_num_col = 7;
  assign cparam_avg_pool_serial_52_act_num_row = 7;
  assign cparam_avg_pool_serial_52_stride_col = 1;
  assign cparam_avg_pool_serial_52_stride_row = 1;
  assign cparam_avg_pool_serial_52_out_num_col = 7;
  assign cparam_avg_pool_serial_52_out_num_row = 7;
  assign cparam_avg_pool_serial_52_pad_col_left = 0;
  assign cparam_avg_pool_serial_52_pad_row_top = 0;
  assign cparam_avg_pool_serial_52_max_col_count = 6;
  assign cparam_avg_pool_serial_52_max_row_count = 6;
  assign cparam_avg_pool_serial_52_max_bat_count = 0;
  assign cparam_avg_pool_serial_52_act_offset_values_0 = 0;
  assign cparam_avg_pool_serial_52_act_row_step = 3584;
  assign cparam_avg_pool_serial_52_act_bat_step = 25088;
  assign cparam_avg_pool_serial_52_act_read_size = 3584;
  assign cparam_avg_pool_serial_52_act_read_block = 512;
  assign cparam_avg_pool_serial_52_out_row_step = 3584;
  assign cparam_avg_pool_serial_52_out_bat_step = 25088;
  assign cparam_avg_pool_serial_52_out_write_size = 3584;
  assign cparam_avg_pool_serial_52_stream_size = 512;
  assign cparam_avg_pool_serial_52_col_select_initval = 0;
  assign cparam_avg_pool_serial_52_stride_col_mod_ksize = 0;
  assign cparam_avg_pool_serial_52_ksize_col_minus_stride_col_mod = 1;
  assign cparam_avg_pool_serial_52_local_pad_offset = 0;
  assign cparam_avg_pool_serial_52_inc_act_laddr = 512;
  assign cparam_avg_pool_serial_52_inc_out_laddr = 512;
  wire [1-1:0] cparam_matmul_55_act_num_col;
  wire [1-1:0] cparam_matmul_55_act_num_row;
  wire [13-1:0] cparam_matmul_55_filter_num_och;
  wire [1-1:0] cparam_matmul_55_bias_scala;
  wire [13-1:0] cparam_matmul_55_bias_num;
  wire [1-1:0] cparam_matmul_55_scale_scala;
  wire [1-1:0] cparam_matmul_55_scale_num;
  wire [1-1:0] cparam_matmul_55_vshamt_mul_scala;
  wire [1-1:0] cparam_matmul_55_vshamt_mul_num;
  wire [1-1:0] cparam_matmul_55_vshamt_sum_scala;
  wire [1-1:0] cparam_matmul_55_vshamt_sum_num;
  wire [1-1:0] cparam_matmul_55_vshamt_out_scala;
  wire [1-1:0] cparam_matmul_55_vshamt_out_num;
  wire [1-1:0] cparam_matmul_55_cshamt_mul_value;
  wire [1-1:0] cparam_matmul_55_cshamt_sum_value;
  wire [5-1:0] cparam_matmul_55_cshamt_out_value;
  wire [1-1:0] cparam_matmul_55_act_func_index;
  wire [1-1:0] cparam_matmul_55_out_num_col;
  wire [1-1:0] cparam_matmul_55_out_num_row;
  wire [1-1:0] cparam_matmul_55_pad_col_left;
  wire [1-1:0] cparam_matmul_55_pad_row_top;
  wire [1-1:0] cparam_matmul_55_max_col_count;
  wire [1-1:0] cparam_matmul_55_max_row_count;
  wire [1-1:0] cparam_matmul_55_max_bat_count;
  wire [12-1:0] cparam_matmul_55_max_och_count;
  wire [6-1:0] cparam_matmul_55_och_count_step;
  wire [1-1:0] cparam_matmul_55_dma_flag_conds_0;
  wire signed [32-1:0] cparam_matmul_55_act_offset_values_0;
  wire [15-1:0] cparam_matmul_55_act_row_step;
  wire [15-1:0] cparam_matmul_55_act_bat_step;
  wire [15-1:0] cparam_matmul_55_act_read_size;
  wire [15-1:0] cparam_matmul_55_act_read_block;
  wire [15-1:0] cparam_matmul_55_act_read_step;
  wire [18-1:0] cparam_matmul_55_filter_base_step;
  wire [18-1:0] cparam_matmul_55_filter_read_size;
  wire [15-1:0] cparam_matmul_55_filter_read_block;
  wire [18-1:0] cparam_matmul_55_filter_read_step;
  wire [1-1:0] cparam_matmul_55_out_offset_values_0;
  wire [13-1:0] cparam_matmul_55_out_col_step;
  wire [13-1:0] cparam_matmul_55_out_row_step;
  wire [13-1:0] cparam_matmul_55_out_bat_step;
  wire [6-1:0] cparam_matmul_55_out_och_step;
  wire [6-1:0] cparam_matmul_55_out_write_size;
  wire [6-1:0] cparam_matmul_55_out_write_size_res;
  wire [1-1:0] cparam_matmul_55_out_write_block;
  wire [1-1:0] cparam_matmul_55_keep_filter;
  wire [1-1:0] cparam_matmul_55_keep_input;
  wire [1-1:0] cparam_matmul_55_data_stationary;
  wire [6-1:0] cparam_matmul_55_stream_num_ops;
  wire [6-1:0] cparam_matmul_55_stream_num_ops_res;
  wire [6-1:0] cparam_matmul_55_stream_num_ops_par;
  wire [6-1:0] cparam_matmul_55_stream_num_ops_res_par;
  wire [15-1:0] cparam_matmul_55_stream_reduce_size;
  wire [15-1:0] cparam_matmul_55_stream_aligned_reduce_size;
  wire [1-1:0] cparam_matmul_55_stream_omit_mask;
  wire [1-1:0] cparam_matmul_55_col_select_initval;
  wire [1-1:0] cparam_matmul_55_stride_col_par_col;
  wire [1-1:0] cparam_matmul_55_stride_row_par_row;
  wire [1-1:0] cparam_matmul_55_stride_col_mod_filter_num;
  wire [1-1:0] cparam_matmul_55_filter_num_col_minus_stride_col_mod;
  wire [1-1:0] cparam_matmul_55_inc_act_laddr_conds_0;
  wire [15-1:0] cparam_matmul_55_inc_act_laddr_small;
  wire [15-1:0] cparam_matmul_55_inc_act_laddr_large;
  wire [13-1:0] cparam_matmul_55_inc_out_laddr_col;
  wire [1-1:0] cparam_matmul_55_stream_act_local_small_offset;
  wire [1-1:0] cparam_matmul_55_stream_act_local_large_offset;
  wire [1-1:0] cparam_matmul_55_stream_act_local_small_flags_0;
  wire [1-1:0] cparam_matmul_55_stream_act_local_large_flags_0;
  wire [1-1:0] cparam_matmul_55_inc_sync_out;
  wire [1-1:0] cparam_matmul_55_inc_sync_out_res;
  reg [2-1:0] matmul_55_control_param_index;
  assign cparam_matmul_55_act_num_col = (matmul_55_control_param_index == 0)? 32'h1 : 
                                        (matmul_55_control_param_index == 1)? 32'h1 : 32'h1;
  assign cparam_matmul_55_act_num_row = (matmul_55_control_param_index == 0)? 32'h1 : 
                                        (matmul_55_control_param_index == 1)? 32'h1 : 32'h1;
  assign cparam_matmul_55_filter_num_och = (matmul_55_control_param_index == 0)? 32'h1000 : 
                                           (matmul_55_control_param_index == 1)? 32'h1000 : 32'h3e8;
  assign cparam_matmul_55_bias_scala = (matmul_55_control_param_index == 0)? 32'h0 : 
                                       (matmul_55_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_matmul_55_bias_num = (matmul_55_control_param_index == 0)? 32'h1000 : 
                                     (matmul_55_control_param_index == 1)? 32'h1000 : 32'h3e8;
  assign cparam_matmul_55_scale_scala = (matmul_55_control_param_index == 0)? 32'h1 : 
                                        (matmul_55_control_param_index == 1)? 32'h1 : 32'h1;
  assign cparam_matmul_55_scale_num = (matmul_55_control_param_index == 0)? 32'h1 : 
                                      (matmul_55_control_param_index == 1)? 32'h1 : 32'h1;
  assign cparam_matmul_55_vshamt_mul_scala = (matmul_55_control_param_index == 0)? 32'h0 : 
                                             (matmul_55_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_matmul_55_vshamt_mul_num = (matmul_55_control_param_index == 0)? 32'h0 : 
                                           (matmul_55_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_matmul_55_vshamt_sum_scala = (matmul_55_control_param_index == 0)? 32'h0 : 
                                             (matmul_55_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_matmul_55_vshamt_sum_num = (matmul_55_control_param_index == 0)? 32'h0 : 
                                           (matmul_55_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_matmul_55_vshamt_out_scala = (matmul_55_control_param_index == 0)? 32'h0 : 
                                             (matmul_55_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_matmul_55_vshamt_out_num = (matmul_55_control_param_index == 0)? 32'h0 : 
                                           (matmul_55_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_matmul_55_cshamt_mul_value = (matmul_55_control_param_index == 0)? 32'h0 : 
                                             (matmul_55_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_matmul_55_cshamt_sum_value = (matmul_55_control_param_index == 0)? 32'h0 : 
                                             (matmul_55_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_matmul_55_cshamt_out_value = (matmul_55_control_param_index == 0)? 32'h11 : 
                                             (matmul_55_control_param_index == 1)? 32'h12 : 32'h12;
  assign cparam_matmul_55_act_func_index = (matmul_55_control_param_index == 0)? 32'h0 : 
                                           (matmul_55_control_param_index == 1)? 32'h0 : 32'h1;
  assign cparam_matmul_55_out_num_col = (matmul_55_control_param_index == 0)? 32'h1 : 
                                        (matmul_55_control_param_index == 1)? 32'h1 : 32'h1;
  assign cparam_matmul_55_out_num_row = (matmul_55_control_param_index == 0)? 32'h1 : 
                                        (matmul_55_control_param_index == 1)? 32'h1 : 32'h1;
  assign cparam_matmul_55_pad_col_left = (matmul_55_control_param_index == 0)? 32'h0 : 
                                         (matmul_55_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_matmul_55_pad_row_top = (matmul_55_control_param_index == 0)? 32'h0 : 
                                        (matmul_55_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_matmul_55_max_col_count = (matmul_55_control_param_index == 0)? 32'h0 : 
                                          (matmul_55_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_matmul_55_max_row_count = (matmul_55_control_param_index == 0)? 32'h0 : 
                                          (matmul_55_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_matmul_55_max_bat_count = (matmul_55_control_param_index == 0)? 32'h0 : 
                                          (matmul_55_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_matmul_55_max_och_count = (matmul_55_control_param_index == 0)? 32'hffc : 
                                          (matmul_55_control_param_index == 1)? 32'hfe0 : 32'h3c8;
  assign cparam_matmul_55_och_count_step = (matmul_55_control_param_index == 0)? 32'h4 : 
                                           (matmul_55_control_param_index == 1)? 32'h20 : 32'h20;
  assign cparam_matmul_55_dma_flag_conds_0 = (matmul_55_control_param_index == 0)? 32'h1 : 
                                             (matmul_55_control_param_index == 1)? 32'h1 : 32'h1;
  assign cparam_matmul_55_act_offset_values_0 = (matmul_55_control_param_index == 0)? 32'h0 : 
                                                (matmul_55_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_matmul_55_act_row_step = (matmul_55_control_param_index == 0)? 32'h6200 : 
                                         (matmul_55_control_param_index == 1)? 32'h1000 : 32'h1000;
  assign cparam_matmul_55_act_bat_step = (matmul_55_control_param_index == 0)? 32'h6200 : 
                                         (matmul_55_control_param_index == 1)? 32'h1000 : 32'h1000;
  assign cparam_matmul_55_act_read_size = (matmul_55_control_param_index == 0)? 32'h6200 : 
                                          (matmul_55_control_param_index == 1)? 32'h1000 : 32'h1000;
  assign cparam_matmul_55_act_read_block = (matmul_55_control_param_index == 0)? 32'h6200 : 
                                           (matmul_55_control_param_index == 1)? 32'h1000 : 32'h1000;
  assign cparam_matmul_55_act_read_step = (matmul_55_control_param_index == 0)? 32'h6200 : 
                                          (matmul_55_control_param_index == 1)? 32'h1000 : 32'h1000;
  assign cparam_matmul_55_filter_base_step = (matmul_55_control_param_index == 0)? 32'h18800 : 
                                             (matmul_55_control_param_index == 1)? 32'h20000 : 32'h20000;
  assign cparam_matmul_55_filter_read_size = (matmul_55_control_param_index == 0)? 32'h18800 : 
                                             (matmul_55_control_param_index == 1)? 32'h20000 : 32'h20000;
  assign cparam_matmul_55_filter_read_block = (matmul_55_control_param_index == 0)? 32'h6200 : 
                                              (matmul_55_control_param_index == 1)? 32'h1000 : 32'h1000;
  assign cparam_matmul_55_filter_read_step = (matmul_55_control_param_index == 0)? 32'h18800 : 
                                             (matmul_55_control_param_index == 1)? 32'h20000 : 32'h20000;
  assign cparam_matmul_55_out_offset_values_0 = (matmul_55_control_param_index == 0)? 32'h0 : 
                                                (matmul_55_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_matmul_55_out_col_step = (matmul_55_control_param_index == 0)? 32'h1000 : 
                                         (matmul_55_control_param_index == 1)? 32'h1000 : 32'h3e8;
  assign cparam_matmul_55_out_row_step = (matmul_55_control_param_index == 0)? 32'h1000 : 
                                         (matmul_55_control_param_index == 1)? 32'h1000 : 32'h3e8;
  assign cparam_matmul_55_out_bat_step = (matmul_55_control_param_index == 0)? 32'h1000 : 
                                         (matmul_55_control_param_index == 1)? 32'h1000 : 32'h3e8;
  assign cparam_matmul_55_out_och_step = (matmul_55_control_param_index == 0)? 32'h4 : 
                                         (matmul_55_control_param_index == 1)? 32'h20 : 32'h20;
  assign cparam_matmul_55_out_write_size = (matmul_55_control_param_index == 0)? 32'h4 : 
                                           (matmul_55_control_param_index == 1)? 32'h20 : 32'h20;
  assign cparam_matmul_55_out_write_size_res = (matmul_55_control_param_index == 0)? 32'h4 : 
                                               (matmul_55_control_param_index == 1)? 32'h20 : 32'h8;
  assign cparam_matmul_55_out_write_block = (matmul_55_control_param_index == 0)? 32'h0 : 
                                            (matmul_55_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_matmul_55_keep_filter = (matmul_55_control_param_index == 0)? 32'h0 : 
                                        (matmul_55_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_matmul_55_keep_input = (matmul_55_control_param_index == 0)? 32'h1 : 
                                       (matmul_55_control_param_index == 1)? 32'h1 : 32'h1;
  assign cparam_matmul_55_data_stationary = (matmul_55_control_param_index == 0)? 32'h0 : 
                                            (matmul_55_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_matmul_55_stream_num_ops = (matmul_55_control_param_index == 0)? 32'h4 : 
                                           (matmul_55_control_param_index == 1)? 32'h20 : 32'h20;
  assign cparam_matmul_55_stream_num_ops_res = (matmul_55_control_param_index == 0)? 32'h4 : 
                                               (matmul_55_control_param_index == 1)? 32'h20 : 32'h8;
  assign cparam_matmul_55_stream_num_ops_par = (matmul_55_control_param_index == 0)? 32'h4 : 
                                               (matmul_55_control_param_index == 1)? 32'h20 : 32'h20;
  assign cparam_matmul_55_stream_num_ops_res_par = (matmul_55_control_param_index == 0)? 32'h4 : 
                                                   (matmul_55_control_param_index == 1)? 32'h20 : 32'h8;
  assign cparam_matmul_55_stream_reduce_size = (matmul_55_control_param_index == 0)? 32'h6200 : 
                                               (matmul_55_control_param_index == 1)? 32'h1000 : 32'h1000;
  assign cparam_matmul_55_stream_aligned_reduce_size = (matmul_55_control_param_index == 0)? 32'h6200 : 
                                                       (matmul_55_control_param_index == 1)? 32'h1000 : 32'h1000;
  assign cparam_matmul_55_stream_omit_mask = (matmul_55_control_param_index == 0)? 32'h0 : 
                                             (matmul_55_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_matmul_55_col_select_initval = (matmul_55_control_param_index == 0)? 32'h0 : 
                                               (matmul_55_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_matmul_55_stride_col_par_col = (matmul_55_control_param_index == 0)? 32'h1 : 
                                               (matmul_55_control_param_index == 1)? 32'h1 : 32'h1;
  assign cparam_matmul_55_stride_row_par_row = (matmul_55_control_param_index == 0)? 32'h1 : 
                                               (matmul_55_control_param_index == 1)? 32'h1 : 32'h1;
  assign cparam_matmul_55_stride_col_mod_filter_num = (matmul_55_control_param_index == 0)? 32'h0 : 
                                                      (matmul_55_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_matmul_55_filter_num_col_minus_stride_col_mod = (matmul_55_control_param_index == 0)? 32'h1 : 
                                                                (matmul_55_control_param_index == 1)? 32'h1 : 32'h1;
  assign cparam_matmul_55_inc_act_laddr_conds_0 = (matmul_55_control_param_index == 0)? 32'h0 : 
                                                  (matmul_55_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_matmul_55_inc_act_laddr_small = (matmul_55_control_param_index == 0)? 32'h6200 : 
                                                (matmul_55_control_param_index == 1)? 32'h1000 : 32'h1000;
  assign cparam_matmul_55_inc_act_laddr_large = (matmul_55_control_param_index == 0)? 32'h6200 : 
                                                (matmul_55_control_param_index == 1)? 32'h1000 : 32'h1000;
  assign cparam_matmul_55_inc_out_laddr_col = (matmul_55_control_param_index == 0)? 32'h1000 : 
                                              (matmul_55_control_param_index == 1)? 32'h1000 : 32'h3e8;
  assign cparam_matmul_55_stream_act_local_small_offset = (matmul_55_control_param_index == 0)? 32'h0 : 
                                                          (matmul_55_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_matmul_55_stream_act_local_large_offset = (matmul_55_control_param_index == 0)? 32'h0 : 
                                                          (matmul_55_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_matmul_55_stream_act_local_small_flags_0 = (matmul_55_control_param_index == 0)? 32'h0 : 
                                                           (matmul_55_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_matmul_55_stream_act_local_large_flags_0 = (matmul_55_control_param_index == 0)? 32'h0 : 
                                                           (matmul_55_control_param_index == 1)? 32'h0 : 32'h0;
  assign cparam_matmul_55_inc_sync_out = (matmul_55_control_param_index == 0)? 32'h1 : 
                                         (matmul_55_control_param_index == 1)? 32'h1 : 32'h1;
  assign cparam_matmul_55_inc_sync_out_res = (matmul_55_control_param_index == 0)? 32'h0 : 
                                             (matmul_55_control_param_index == 1)? 32'h0 : 32'h0;
  reg _acc_0_stream_ivalid;
  wire _acc_0_stream_oready;
  wire _acc_0_stream_internal_oready;
  assign _acc_0_stream_internal_oready = 1;
  reg [32-1:0] _acc_0_fsm;
  localparam _acc_0_fsm_init = 0;
  wire _acc_0_run_flag;
  assign _acc_0_run_flag = 0;
  reg _acc_0_source_start;
  wire _acc_0_source_stop;
  reg _acc_0_source_busy;
  wire _acc_0_sink_start;
  wire _acc_0_sink_stop;
  wire _acc_0_sink_busy;
  wire _acc_0_busy;
  reg _acc_0_busy_reg;
  wire _acc_0_is_root;
  reg _acc_0_x_idle;
  reg [33-1:0] _acc_0_x_source_count;
  reg [5-1:0] _acc_0_x_source_mode;
  reg [16-1:0] _acc_0_x_source_generator_id;
  reg [32-1:0] _acc_0_x_source_offset;
  reg [33-1:0] _acc_0_x_source_size;
  reg [32-1:0] _acc_0_x_source_stride;
  reg [32-1:0] _acc_0_x_source_offset_buf;
  reg [33-1:0] _acc_0_x_source_size_buf;
  reg [32-1:0] _acc_0_x_source_stride_buf;
  reg [8-1:0] _acc_0_x_source_sel;
  reg [32-1:0] _acc_0_x_source_ram_raddr;
  reg _acc_0_x_source_ram_renable;
  wire [32-1:0] _acc_0_x_source_ram_rdata;
  reg _acc_0_x_source_fifo_deq;
  wire [32-1:0] _acc_0_x_source_fifo_rdata;
  reg [32-1:0] _acc_0_x_source_empty_data;
  reg _acc_0_rshift_idle;
  reg [33-1:0] _acc_0_rshift_source_count;
  reg [5-1:0] _acc_0_rshift_source_mode;
  reg [16-1:0] _acc_0_rshift_source_generator_id;
  reg [32-1:0] _acc_0_rshift_source_offset;
  reg [33-1:0] _acc_0_rshift_source_size;
  reg [32-1:0] _acc_0_rshift_source_stride;
  reg [32-1:0] _acc_0_rshift_source_offset_buf;
  reg [33-1:0] _acc_0_rshift_source_size_buf;
  reg [32-1:0] _acc_0_rshift_source_stride_buf;
  reg [8-1:0] _acc_0_rshift_source_sel;
  reg [32-1:0] _acc_0_rshift_source_ram_raddr;
  reg _acc_0_rshift_source_ram_renable;
  wire [32-1:0] _acc_0_rshift_source_ram_rdata;
  reg _acc_0_rshift_source_fifo_deq;
  wire [32-1:0] _acc_0_rshift_source_fifo_rdata;
  reg [32-1:0] _acc_0_rshift_source_empty_data;
  reg [32-1:0] _acc_0_size_next_parameter_data;
  reg [33-1:0] _acc_0_sum_sink_count;
  reg [5-1:0] _acc_0_sum_sink_mode;
  reg [16-1:0] _acc_0_sum_sink_generator_id;
  reg [32-1:0] _acc_0_sum_sink_offset;
  reg [33-1:0] _acc_0_sum_sink_size;
  reg [32-1:0] _acc_0_sum_sink_stride;
  reg [32-1:0] _acc_0_sum_sink_offset_buf;
  reg [33-1:0] _acc_0_sum_sink_size_buf;
  reg [32-1:0] _acc_0_sum_sink_stride_buf;
  reg [8-1:0] _acc_0_sum_sink_sel;
  reg [32-1:0] _acc_0_sum_sink_waddr;
  reg _acc_0_sum_sink_wenable;
  reg [32-1:0] _acc_0_sum_sink_wdata;
  reg _acc_0_sum_sink_fifo_enq;
  reg [32-1:0] _acc_0_sum_sink_fifo_wdata;
  reg [32-1:0] _acc_0_sum_sink_immediate;
  reg [33-1:0] _acc_0_valid_sink_count;
  reg [5-1:0] _acc_0_valid_sink_mode;
  reg [16-1:0] _acc_0_valid_sink_generator_id;
  reg [32-1:0] _acc_0_valid_sink_offset;
  reg [33-1:0] _acc_0_valid_sink_size;
  reg [32-1:0] _acc_0_valid_sink_stride;
  reg [32-1:0] _acc_0_valid_sink_offset_buf;
  reg [33-1:0] _acc_0_valid_sink_size_buf;
  reg [32-1:0] _acc_0_valid_sink_stride_buf;
  reg [8-1:0] _acc_0_valid_sink_sel;
  reg [32-1:0] _acc_0_valid_sink_waddr;
  reg _acc_0_valid_sink_wenable;
  reg [1-1:0] _acc_0_valid_sink_wdata;
  reg _acc_0_valid_sink_fifo_enq;
  reg [1-1:0] _acc_0_valid_sink_fifo_wdata;
  reg [1-1:0] _acc_0_valid_sink_immediate;
  reg _acc_1_stream_ivalid;
  wire _acc_1_stream_oready;
  wire _acc_1_stream_internal_oready;
  assign _acc_1_stream_internal_oready = 1;
  reg [32-1:0] _acc_1_fsm;
  localparam _acc_1_fsm_init = 0;
  wire _acc_1_run_flag;
  assign _acc_1_run_flag = 0;
  reg _acc_1_source_start;
  wire _acc_1_source_stop;
  reg _acc_1_source_busy;
  wire _acc_1_sink_start;
  wire _acc_1_sink_stop;
  wire _acc_1_sink_busy;
  wire _acc_1_busy;
  reg _acc_1_busy_reg;
  wire _acc_1_is_root;
  reg _acc_1_x_idle;
  reg [33-1:0] _acc_1_x_source_count;
  reg [5-1:0] _acc_1_x_source_mode;
  reg [16-1:0] _acc_1_x_source_generator_id;
  reg [32-1:0] _acc_1_x_source_offset;
  reg [33-1:0] _acc_1_x_source_size;
  reg [32-1:0] _acc_1_x_source_stride;
  reg [32-1:0] _acc_1_x_source_offset_buf;
  reg [33-1:0] _acc_1_x_source_size_buf;
  reg [32-1:0] _acc_1_x_source_stride_buf;
  reg [8-1:0] _acc_1_x_source_sel;
  reg [32-1:0] _acc_1_x_source_ram_raddr;
  reg _acc_1_x_source_ram_renable;
  wire [32-1:0] _acc_1_x_source_ram_rdata;
  reg _acc_1_x_source_fifo_deq;
  wire [32-1:0] _acc_1_x_source_fifo_rdata;
  reg [32-1:0] _acc_1_x_source_empty_data;
  reg _acc_1_rshift_idle;
  reg [33-1:0] _acc_1_rshift_source_count;
  reg [5-1:0] _acc_1_rshift_source_mode;
  reg [16-1:0] _acc_1_rshift_source_generator_id;
  reg [32-1:0] _acc_1_rshift_source_offset;
  reg [33-1:0] _acc_1_rshift_source_size;
  reg [32-1:0] _acc_1_rshift_source_stride;
  reg [32-1:0] _acc_1_rshift_source_offset_buf;
  reg [33-1:0] _acc_1_rshift_source_size_buf;
  reg [32-1:0] _acc_1_rshift_source_stride_buf;
  reg [8-1:0] _acc_1_rshift_source_sel;
  reg [32-1:0] _acc_1_rshift_source_ram_raddr;
  reg _acc_1_rshift_source_ram_renable;
  wire [32-1:0] _acc_1_rshift_source_ram_rdata;
  reg _acc_1_rshift_source_fifo_deq;
  wire [32-1:0] _acc_1_rshift_source_fifo_rdata;
  reg [32-1:0] _acc_1_rshift_source_empty_data;
  reg [32-1:0] _acc_1_size_next_parameter_data;
  reg [33-1:0] _acc_1_sum_sink_count;
  reg [5-1:0] _acc_1_sum_sink_mode;
  reg [16-1:0] _acc_1_sum_sink_generator_id;
  reg [32-1:0] _acc_1_sum_sink_offset;
  reg [33-1:0] _acc_1_sum_sink_size;
  reg [32-1:0] _acc_1_sum_sink_stride;
  reg [32-1:0] _acc_1_sum_sink_offset_buf;
  reg [33-1:0] _acc_1_sum_sink_size_buf;
  reg [32-1:0] _acc_1_sum_sink_stride_buf;
  reg [8-1:0] _acc_1_sum_sink_sel;
  reg [32-1:0] _acc_1_sum_sink_waddr;
  reg _acc_1_sum_sink_wenable;
  reg [32-1:0] _acc_1_sum_sink_wdata;
  reg _acc_1_sum_sink_fifo_enq;
  reg [32-1:0] _acc_1_sum_sink_fifo_wdata;
  reg [32-1:0] _acc_1_sum_sink_immediate;
  reg [33-1:0] _acc_1_valid_sink_count;
  reg [5-1:0] _acc_1_valid_sink_mode;
  reg [16-1:0] _acc_1_valid_sink_generator_id;
  reg [32-1:0] _acc_1_valid_sink_offset;
  reg [33-1:0] _acc_1_valid_sink_size;
  reg [32-1:0] _acc_1_valid_sink_stride;
  reg [32-1:0] _acc_1_valid_sink_offset_buf;
  reg [33-1:0] _acc_1_valid_sink_size_buf;
  reg [32-1:0] _acc_1_valid_sink_stride_buf;
  reg [8-1:0] _acc_1_valid_sink_sel;
  reg [32-1:0] _acc_1_valid_sink_waddr;
  reg _acc_1_valid_sink_wenable;
  reg [1-1:0] _acc_1_valid_sink_wdata;
  reg _acc_1_valid_sink_fifo_enq;
  reg [1-1:0] _acc_1_valid_sink_fifo_wdata;
  reg [1-1:0] _acc_1_valid_sink_immediate;
  reg _add_tree_2_stream_ivalid;
  wire _add_tree_2_stream_oready;
  wire _add_tree_2_stream_internal_oready;
  assign _add_tree_2_stream_internal_oready = 1;
  reg [32-1:0] _add_tree_2_fsm;
  localparam _add_tree_2_fsm_init = 0;
  wire _add_tree_2_run_flag;
  assign _add_tree_2_run_flag = 0;
  reg _add_tree_2_source_start;
  wire _add_tree_2_source_stop;
  reg _add_tree_2_source_busy;
  wire _add_tree_2_sink_start;
  wire _add_tree_2_sink_stop;
  wire _add_tree_2_sink_busy;
  wire _add_tree_2_busy;
  reg _add_tree_2_busy_reg;
  wire _add_tree_2_is_root;
  reg _add_tree_2_var0_idle;
  reg [33-1:0] _add_tree_2_var0_source_count;
  reg [5-1:0] _add_tree_2_var0_source_mode;
  reg [16-1:0] _add_tree_2_var0_source_generator_id;
  reg [32-1:0] _add_tree_2_var0_source_offset;
  reg [33-1:0] _add_tree_2_var0_source_size;
  reg [32-1:0] _add_tree_2_var0_source_stride;
  reg [32-1:0] _add_tree_2_var0_source_offset_buf;
  reg [33-1:0] _add_tree_2_var0_source_size_buf;
  reg [32-1:0] _add_tree_2_var0_source_stride_buf;
  reg [8-1:0] _add_tree_2_var0_source_sel;
  reg [32-1:0] _add_tree_2_var0_source_ram_raddr;
  reg _add_tree_2_var0_source_ram_renable;
  wire [32-1:0] _add_tree_2_var0_source_ram_rdata;
  reg _add_tree_2_var0_source_fifo_deq;
  wire [32-1:0] _add_tree_2_var0_source_fifo_rdata;
  reg [32-1:0] _add_tree_2_var0_source_empty_data;
  reg [33-1:0] _add_tree_2_sum_sink_count;
  reg [5-1:0] _add_tree_2_sum_sink_mode;
  reg [16-1:0] _add_tree_2_sum_sink_generator_id;
  reg [32-1:0] _add_tree_2_sum_sink_offset;
  reg [33-1:0] _add_tree_2_sum_sink_size;
  reg [32-1:0] _add_tree_2_sum_sink_stride;
  reg [32-1:0] _add_tree_2_sum_sink_offset_buf;
  reg [33-1:0] _add_tree_2_sum_sink_size_buf;
  reg [32-1:0] _add_tree_2_sum_sink_stride_buf;
  reg [8-1:0] _add_tree_2_sum_sink_sel;
  reg [32-1:0] _add_tree_2_sum_sink_waddr;
  reg _add_tree_2_sum_sink_wenable;
  reg [32-1:0] _add_tree_2_sum_sink_wdata;
  reg _add_tree_2_sum_sink_fifo_enq;
  reg [32-1:0] _add_tree_2_sum_sink_fifo_wdata;
  reg [32-1:0] _add_tree_2_sum_sink_immediate;
  reg _add_tree_3_stream_ivalid;
  wire _add_tree_3_stream_oready;
  wire _add_tree_3_stream_internal_oready;
  assign _add_tree_3_stream_internal_oready = 1;
  reg [32-1:0] _add_tree_3_fsm;
  localparam _add_tree_3_fsm_init = 0;
  wire _add_tree_3_run_flag;
  assign _add_tree_3_run_flag = 0;
  reg _add_tree_3_source_start;
  wire _add_tree_3_source_stop;
  reg _add_tree_3_source_busy;
  wire _add_tree_3_sink_start;
  wire _add_tree_3_sink_stop;
  wire _add_tree_3_sink_busy;
  wire _add_tree_3_busy;
  reg _add_tree_3_busy_reg;
  wire _add_tree_3_is_root;
  reg _add_tree_3_var0_idle;
  reg [33-1:0] _add_tree_3_var0_source_count;
  reg [5-1:0] _add_tree_3_var0_source_mode;
  reg [16-1:0] _add_tree_3_var0_source_generator_id;
  reg [32-1:0] _add_tree_3_var0_source_offset;
  reg [33-1:0] _add_tree_3_var0_source_size;
  reg [32-1:0] _add_tree_3_var0_source_stride;
  reg [32-1:0] _add_tree_3_var0_source_offset_buf;
  reg [33-1:0] _add_tree_3_var0_source_size_buf;
  reg [32-1:0] _add_tree_3_var0_source_stride_buf;
  reg [8-1:0] _add_tree_3_var0_source_sel;
  reg [32-1:0] _add_tree_3_var0_source_ram_raddr;
  reg _add_tree_3_var0_source_ram_renable;
  wire [32-1:0] _add_tree_3_var0_source_ram_rdata;
  reg _add_tree_3_var0_source_fifo_deq;
  wire [32-1:0] _add_tree_3_var0_source_fifo_rdata;
  reg [32-1:0] _add_tree_3_var0_source_empty_data;
  reg _add_tree_3_var1_idle;
  reg [33-1:0] _add_tree_3_var1_source_count;
  reg [5-1:0] _add_tree_3_var1_source_mode;
  reg [16-1:0] _add_tree_3_var1_source_generator_id;
  reg [32-1:0] _add_tree_3_var1_source_offset;
  reg [33-1:0] _add_tree_3_var1_source_size;
  reg [32-1:0] _add_tree_3_var1_source_stride;
  reg [32-1:0] _add_tree_3_var1_source_offset_buf;
  reg [33-1:0] _add_tree_3_var1_source_size_buf;
  reg [32-1:0] _add_tree_3_var1_source_stride_buf;
  reg [8-1:0] _add_tree_3_var1_source_sel;
  reg [32-1:0] _add_tree_3_var1_source_ram_raddr;
  reg _add_tree_3_var1_source_ram_renable;
  wire [32-1:0] _add_tree_3_var1_source_ram_rdata;
  reg _add_tree_3_var1_source_fifo_deq;
  wire [32-1:0] _add_tree_3_var1_source_fifo_rdata;
  reg [32-1:0] _add_tree_3_var1_source_empty_data;
  reg _add_tree_3_var2_idle;
  reg [33-1:0] _add_tree_3_var2_source_count;
  reg [5-1:0] _add_tree_3_var2_source_mode;
  reg [16-1:0] _add_tree_3_var2_source_generator_id;
  reg [32-1:0] _add_tree_3_var2_source_offset;
  reg [33-1:0] _add_tree_3_var2_source_size;
  reg [32-1:0] _add_tree_3_var2_source_stride;
  reg [32-1:0] _add_tree_3_var2_source_offset_buf;
  reg [33-1:0] _add_tree_3_var2_source_size_buf;
  reg [32-1:0] _add_tree_3_var2_source_stride_buf;
  reg [8-1:0] _add_tree_3_var2_source_sel;
  reg [32-1:0] _add_tree_3_var2_source_ram_raddr;
  reg _add_tree_3_var2_source_ram_renable;
  wire [32-1:0] _add_tree_3_var2_source_ram_rdata;
  reg _add_tree_3_var2_source_fifo_deq;
  wire [32-1:0] _add_tree_3_var2_source_fifo_rdata;
  reg [32-1:0] _add_tree_3_var2_source_empty_data;
  reg _add_tree_3_var3_idle;
  reg [33-1:0] _add_tree_3_var3_source_count;
  reg [5-1:0] _add_tree_3_var3_source_mode;
  reg [16-1:0] _add_tree_3_var3_source_generator_id;
  reg [32-1:0] _add_tree_3_var3_source_offset;
  reg [33-1:0] _add_tree_3_var3_source_size;
  reg [32-1:0] _add_tree_3_var3_source_stride;
  reg [32-1:0] _add_tree_3_var3_source_offset_buf;
  reg [33-1:0] _add_tree_3_var3_source_size_buf;
  reg [32-1:0] _add_tree_3_var3_source_stride_buf;
  reg [8-1:0] _add_tree_3_var3_source_sel;
  reg [32-1:0] _add_tree_3_var3_source_ram_raddr;
  reg _add_tree_3_var3_source_ram_renable;
  wire [32-1:0] _add_tree_3_var3_source_ram_rdata;
  reg _add_tree_3_var3_source_fifo_deq;
  wire [32-1:0] _add_tree_3_var3_source_fifo_rdata;
  reg [32-1:0] _add_tree_3_var3_source_empty_data;
  reg _add_tree_3_var4_idle;
  reg [33-1:0] _add_tree_3_var4_source_count;
  reg [5-1:0] _add_tree_3_var4_source_mode;
  reg [16-1:0] _add_tree_3_var4_source_generator_id;
  reg [32-1:0] _add_tree_3_var4_source_offset;
  reg [33-1:0] _add_tree_3_var4_source_size;
  reg [32-1:0] _add_tree_3_var4_source_stride;
  reg [32-1:0] _add_tree_3_var4_source_offset_buf;
  reg [33-1:0] _add_tree_3_var4_source_size_buf;
  reg [32-1:0] _add_tree_3_var4_source_stride_buf;
  reg [8-1:0] _add_tree_3_var4_source_sel;
  reg [32-1:0] _add_tree_3_var4_source_ram_raddr;
  reg _add_tree_3_var4_source_ram_renable;
  wire [32-1:0] _add_tree_3_var4_source_ram_rdata;
  reg _add_tree_3_var4_source_fifo_deq;
  wire [32-1:0] _add_tree_3_var4_source_fifo_rdata;
  reg [32-1:0] _add_tree_3_var4_source_empty_data;
  reg _add_tree_3_var5_idle;
  reg [33-1:0] _add_tree_3_var5_source_count;
  reg [5-1:0] _add_tree_3_var5_source_mode;
  reg [16-1:0] _add_tree_3_var5_source_generator_id;
  reg [32-1:0] _add_tree_3_var5_source_offset;
  reg [33-1:0] _add_tree_3_var5_source_size;
  reg [32-1:0] _add_tree_3_var5_source_stride;
  reg [32-1:0] _add_tree_3_var5_source_offset_buf;
  reg [33-1:0] _add_tree_3_var5_source_size_buf;
  reg [32-1:0] _add_tree_3_var5_source_stride_buf;
  reg [8-1:0] _add_tree_3_var5_source_sel;
  reg [32-1:0] _add_tree_3_var5_source_ram_raddr;
  reg _add_tree_3_var5_source_ram_renable;
  wire [32-1:0] _add_tree_3_var5_source_ram_rdata;
  reg _add_tree_3_var5_source_fifo_deq;
  wire [32-1:0] _add_tree_3_var5_source_fifo_rdata;
  reg [32-1:0] _add_tree_3_var5_source_empty_data;
  reg _add_tree_3_var6_idle;
  reg [33-1:0] _add_tree_3_var6_source_count;
  reg [5-1:0] _add_tree_3_var6_source_mode;
  reg [16-1:0] _add_tree_3_var6_source_generator_id;
  reg [32-1:0] _add_tree_3_var6_source_offset;
  reg [33-1:0] _add_tree_3_var6_source_size;
  reg [32-1:0] _add_tree_3_var6_source_stride;
  reg [32-1:0] _add_tree_3_var6_source_offset_buf;
  reg [33-1:0] _add_tree_3_var6_source_size_buf;
  reg [32-1:0] _add_tree_3_var6_source_stride_buf;
  reg [8-1:0] _add_tree_3_var6_source_sel;
  reg [32-1:0] _add_tree_3_var6_source_ram_raddr;
  reg _add_tree_3_var6_source_ram_renable;
  wire [32-1:0] _add_tree_3_var6_source_ram_rdata;
  reg _add_tree_3_var6_source_fifo_deq;
  wire [32-1:0] _add_tree_3_var6_source_fifo_rdata;
  reg [32-1:0] _add_tree_3_var6_source_empty_data;
  reg _add_tree_3_var7_idle;
  reg [33-1:0] _add_tree_3_var7_source_count;
  reg [5-1:0] _add_tree_3_var7_source_mode;
  reg [16-1:0] _add_tree_3_var7_source_generator_id;
  reg [32-1:0] _add_tree_3_var7_source_offset;
  reg [33-1:0] _add_tree_3_var7_source_size;
  reg [32-1:0] _add_tree_3_var7_source_stride;
  reg [32-1:0] _add_tree_3_var7_source_offset_buf;
  reg [33-1:0] _add_tree_3_var7_source_size_buf;
  reg [32-1:0] _add_tree_3_var7_source_stride_buf;
  reg [8-1:0] _add_tree_3_var7_source_sel;
  reg [32-1:0] _add_tree_3_var7_source_ram_raddr;
  reg _add_tree_3_var7_source_ram_renable;
  wire [32-1:0] _add_tree_3_var7_source_ram_rdata;
  reg _add_tree_3_var7_source_fifo_deq;
  wire [32-1:0] _add_tree_3_var7_source_fifo_rdata;
  reg [32-1:0] _add_tree_3_var7_source_empty_data;
  reg _add_tree_3_var8_idle;
  reg [33-1:0] _add_tree_3_var8_source_count;
  reg [5-1:0] _add_tree_3_var8_source_mode;
  reg [16-1:0] _add_tree_3_var8_source_generator_id;
  reg [32-1:0] _add_tree_3_var8_source_offset;
  reg [33-1:0] _add_tree_3_var8_source_size;
  reg [32-1:0] _add_tree_3_var8_source_stride;
  reg [32-1:0] _add_tree_3_var8_source_offset_buf;
  reg [33-1:0] _add_tree_3_var8_source_size_buf;
  reg [32-1:0] _add_tree_3_var8_source_stride_buf;
  reg [8-1:0] _add_tree_3_var8_source_sel;
  reg [32-1:0] _add_tree_3_var8_source_ram_raddr;
  reg _add_tree_3_var8_source_ram_renable;
  wire [32-1:0] _add_tree_3_var8_source_ram_rdata;
  reg _add_tree_3_var8_source_fifo_deq;
  wire [32-1:0] _add_tree_3_var8_source_fifo_rdata;
  reg [32-1:0] _add_tree_3_var8_source_empty_data;
  reg [33-1:0] _add_tree_3_sum_sink_count;
  reg [5-1:0] _add_tree_3_sum_sink_mode;
  reg [16-1:0] _add_tree_3_sum_sink_generator_id;
  reg [32-1:0] _add_tree_3_sum_sink_offset;
  reg [33-1:0] _add_tree_3_sum_sink_size;
  reg [32-1:0] _add_tree_3_sum_sink_stride;
  reg [32-1:0] _add_tree_3_sum_sink_offset_buf;
  reg [33-1:0] _add_tree_3_sum_sink_size_buf;
  reg [32-1:0] _add_tree_3_sum_sink_stride_buf;
  reg [8-1:0] _add_tree_3_sum_sink_sel;
  reg [32-1:0] _add_tree_3_sum_sink_waddr;
  reg _add_tree_3_sum_sink_wenable;
  reg [32-1:0] _add_tree_3_sum_sink_wdata;
  reg _add_tree_3_sum_sink_fifo_enq;
  reg [32-1:0] _add_tree_3_sum_sink_fifo_wdata;
  reg [32-1:0] _add_tree_3_sum_sink_immediate;
  reg _mul_rshift_round_clip_4_stream_ivalid;
  wire _mul_rshift_round_clip_4_stream_oready;
  wire _mul_rshift_round_clip_4_stream_internal_oready;
  assign _mul_rshift_round_clip_4_stream_internal_oready = 1;
  reg [32-1:0] _mul_rshift_round_clip_4_fsm;
  localparam _mul_rshift_round_clip_4_fsm_init = 0;
  wire _mul_rshift_round_clip_4_run_flag;
  assign _mul_rshift_round_clip_4_run_flag = 0;
  reg _mul_rshift_round_clip_4_source_start;
  wire _mul_rshift_round_clip_4_source_stop;
  reg _mul_rshift_round_clip_4_source_busy;
  wire _mul_rshift_round_clip_4_sink_start;
  wire _mul_rshift_round_clip_4_sink_stop;
  wire _mul_rshift_round_clip_4_sink_busy;
  wire _mul_rshift_round_clip_4_busy;
  reg _mul_rshift_round_clip_4_busy_reg;
  wire _mul_rshift_round_clip_4_is_root;
  reg _mul_rshift_round_clip_4_x_idle;
  reg [33-1:0] _mul_rshift_round_clip_4_x_source_count;
  reg [5-1:0] _mul_rshift_round_clip_4_x_source_mode;
  reg [16-1:0] _mul_rshift_round_clip_4_x_source_generator_id;
  reg [32-1:0] _mul_rshift_round_clip_4_x_source_offset;
  reg [33-1:0] _mul_rshift_round_clip_4_x_source_size;
  reg [32-1:0] _mul_rshift_round_clip_4_x_source_stride;
  reg [32-1:0] _mul_rshift_round_clip_4_x_source_offset_buf;
  reg [33-1:0] _mul_rshift_round_clip_4_x_source_size_buf;
  reg [32-1:0] _mul_rshift_round_clip_4_x_source_stride_buf;
  reg [8-1:0] _mul_rshift_round_clip_4_x_source_sel;
  reg [32-1:0] _mul_rshift_round_clip_4_x_source_ram_raddr;
  reg _mul_rshift_round_clip_4_x_source_ram_renable;
  wire [32-1:0] _mul_rshift_round_clip_4_x_source_ram_rdata;
  reg _mul_rshift_round_clip_4_x_source_fifo_deq;
  wire [32-1:0] _mul_rshift_round_clip_4_x_source_fifo_rdata;
  reg [32-1:0] _mul_rshift_round_clip_4_x_source_empty_data;
  reg _mul_rshift_round_clip_4_y_idle;
  reg [33-1:0] _mul_rshift_round_clip_4_y_source_count;
  reg [5-1:0] _mul_rshift_round_clip_4_y_source_mode;
  reg [16-1:0] _mul_rshift_round_clip_4_y_source_generator_id;
  reg [32-1:0] _mul_rshift_round_clip_4_y_source_offset;
  reg [33-1:0] _mul_rshift_round_clip_4_y_source_size;
  reg [32-1:0] _mul_rshift_round_clip_4_y_source_stride;
  reg [32-1:0] _mul_rshift_round_clip_4_y_source_offset_buf;
  reg [33-1:0] _mul_rshift_round_clip_4_y_source_size_buf;
  reg [32-1:0] _mul_rshift_round_clip_4_y_source_stride_buf;
  reg [8-1:0] _mul_rshift_round_clip_4_y_source_sel;
  reg [32-1:0] _mul_rshift_round_clip_4_y_source_ram_raddr;
  reg _mul_rshift_round_clip_4_y_source_ram_renable;
  wire [8-1:0] _mul_rshift_round_clip_4_y_source_ram_rdata;
  reg _mul_rshift_round_clip_4_y_source_fifo_deq;
  wire [8-1:0] _mul_rshift_round_clip_4_y_source_fifo_rdata;
  reg [8-1:0] _mul_rshift_round_clip_4_y_source_empty_data;
  reg _mul_rshift_round_clip_4_rshift_idle;
  reg [33-1:0] _mul_rshift_round_clip_4_rshift_source_count;
  reg [5-1:0] _mul_rshift_round_clip_4_rshift_source_mode;
  reg [16-1:0] _mul_rshift_round_clip_4_rshift_source_generator_id;
  reg [32-1:0] _mul_rshift_round_clip_4_rshift_source_offset;
  reg [33-1:0] _mul_rshift_round_clip_4_rshift_source_size;
  reg [32-1:0] _mul_rshift_round_clip_4_rshift_source_stride;
  reg [32-1:0] _mul_rshift_round_clip_4_rshift_source_offset_buf;
  reg [33-1:0] _mul_rshift_round_clip_4_rshift_source_size_buf;
  reg [32-1:0] _mul_rshift_round_clip_4_rshift_source_stride_buf;
  reg [8-1:0] _mul_rshift_round_clip_4_rshift_source_sel;
  reg [32-1:0] _mul_rshift_round_clip_4_rshift_source_ram_raddr;
  reg _mul_rshift_round_clip_4_rshift_source_ram_renable;
  wire [32-1:0] _mul_rshift_round_clip_4_rshift_source_ram_rdata;
  reg _mul_rshift_round_clip_4_rshift_source_fifo_deq;
  wire [32-1:0] _mul_rshift_round_clip_4_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_rshift_round_clip_4_rshift_source_empty_data;
  reg [33-1:0] _mul_rshift_round_clip_4_z_sink_count;
  reg [5-1:0] _mul_rshift_round_clip_4_z_sink_mode;
  reg [16-1:0] _mul_rshift_round_clip_4_z_sink_generator_id;
  reg [32-1:0] _mul_rshift_round_clip_4_z_sink_offset;
  reg [33-1:0] _mul_rshift_round_clip_4_z_sink_size;
  reg [32-1:0] _mul_rshift_round_clip_4_z_sink_stride;
  reg [32-1:0] _mul_rshift_round_clip_4_z_sink_offset_buf;
  reg [33-1:0] _mul_rshift_round_clip_4_z_sink_size_buf;
  reg [32-1:0] _mul_rshift_round_clip_4_z_sink_stride_buf;
  reg [8-1:0] _mul_rshift_round_clip_4_z_sink_sel;
  reg [32-1:0] _mul_rshift_round_clip_4_z_sink_waddr;
  reg _mul_rshift_round_clip_4_z_sink_wenable;
  reg [8-1:0] _mul_rshift_round_clip_4_z_sink_wdata;
  reg _mul_rshift_round_clip_4_z_sink_fifo_enq;
  reg [8-1:0] _mul_rshift_round_clip_4_z_sink_fifo_wdata;
  reg [8-1:0] _mul_rshift_round_clip_4_z_sink_immediate;
  reg _mul_5_stream_ivalid;
  wire _mul_5_stream_oready;
  wire _mul_5_stream_internal_oready;
  assign _mul_5_stream_internal_oready = 1;
  reg [32-1:0] _mul_5_fsm;
  localparam _mul_5_fsm_init = 0;
  wire _mul_5_run_flag;
  assign _mul_5_run_flag = 0;
  reg _mul_5_source_start;
  wire _mul_5_source_stop;
  reg _mul_5_source_busy;
  wire _mul_5_sink_start;
  wire _mul_5_sink_stop;
  wire _mul_5_sink_busy;
  wire _mul_5_busy;
  reg _mul_5_busy_reg;
  wire _mul_5_is_root;
  reg _mul_5_x_idle;
  reg [33-1:0] _mul_5_x_source_count;
  reg [5-1:0] _mul_5_x_source_mode;
  reg [16-1:0] _mul_5_x_source_generator_id;
  reg [32-1:0] _mul_5_x_source_offset;
  reg [33-1:0] _mul_5_x_source_size;
  reg [32-1:0] _mul_5_x_source_stride;
  reg [32-1:0] _mul_5_x_source_offset_buf;
  reg [33-1:0] _mul_5_x_source_size_buf;
  reg [32-1:0] _mul_5_x_source_stride_buf;
  reg [8-1:0] _mul_5_x_source_sel;
  reg [32-1:0] _mul_5_x_source_ram_raddr;
  reg _mul_5_x_source_ram_renable;
  wire [8-1:0] _mul_5_x_source_ram_rdata;
  reg _mul_5_x_source_fifo_deq;
  wire [8-1:0] _mul_5_x_source_fifo_rdata;
  reg [8-1:0] _mul_5_x_source_empty_data;
  reg _mul_5_y_idle;
  reg [33-1:0] _mul_5_y_source_count;
  reg [5-1:0] _mul_5_y_source_mode;
  reg [16-1:0] _mul_5_y_source_generator_id;
  reg [32-1:0] _mul_5_y_source_offset;
  reg [33-1:0] _mul_5_y_source_size;
  reg [32-1:0] _mul_5_y_source_stride;
  reg [32-1:0] _mul_5_y_source_offset_buf;
  reg [33-1:0] _mul_5_y_source_size_buf;
  reg [32-1:0] _mul_5_y_source_stride_buf;
  reg [8-1:0] _mul_5_y_source_sel;
  reg [32-1:0] _mul_5_y_source_ram_raddr;
  reg _mul_5_y_source_ram_renable;
  wire [8-1:0] _mul_5_y_source_ram_rdata;
  reg _mul_5_y_source_fifo_deq;
  wire [8-1:0] _mul_5_y_source_fifo_rdata;
  reg [8-1:0] _mul_5_y_source_empty_data;
  reg _mul_5_rshift_idle;
  reg [33-1:0] _mul_5_rshift_source_count;
  reg [5-1:0] _mul_5_rshift_source_mode;
  reg [16-1:0] _mul_5_rshift_source_generator_id;
  reg [32-1:0] _mul_5_rshift_source_offset;
  reg [33-1:0] _mul_5_rshift_source_size;
  reg [32-1:0] _mul_5_rshift_source_stride;
  reg [32-1:0] _mul_5_rshift_source_offset_buf;
  reg [33-1:0] _mul_5_rshift_source_size_buf;
  reg [32-1:0] _mul_5_rshift_source_stride_buf;
  reg [8-1:0] _mul_5_rshift_source_sel;
  reg [32-1:0] _mul_5_rshift_source_ram_raddr;
  reg _mul_5_rshift_source_ram_renable;
  wire [32-1:0] _mul_5_rshift_source_ram_rdata;
  reg _mul_5_rshift_source_fifo_deq;
  wire [32-1:0] _mul_5_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_5_rshift_source_empty_data;
  reg [33-1:0] _mul_5_z_sink_count;
  reg [5-1:0] _mul_5_z_sink_mode;
  reg [16-1:0] _mul_5_z_sink_generator_id;
  reg [32-1:0] _mul_5_z_sink_offset;
  reg [33-1:0] _mul_5_z_sink_size;
  reg [32-1:0] _mul_5_z_sink_stride;
  reg [32-1:0] _mul_5_z_sink_offset_buf;
  reg [33-1:0] _mul_5_z_sink_size_buf;
  reg [32-1:0] _mul_5_z_sink_stride_buf;
  reg [8-1:0] _mul_5_z_sink_sel;
  reg [32-1:0] _mul_5_z_sink_waddr;
  reg _mul_5_z_sink_wenable;
  reg [16-1:0] _mul_5_z_sink_wdata;
  reg _mul_5_z_sink_fifo_enq;
  reg [16-1:0] _mul_5_z_sink_fifo_wdata;
  reg [16-1:0] _mul_5_z_sink_immediate;
  reg _mul_6_stream_ivalid;
  wire _mul_6_stream_oready;
  wire _mul_6_stream_internal_oready;
  assign _mul_6_stream_internal_oready = 1;
  reg [32-1:0] _mul_6_fsm;
  localparam _mul_6_fsm_init = 0;
  wire _mul_6_run_flag;
  assign _mul_6_run_flag = 0;
  reg _mul_6_source_start;
  wire _mul_6_source_stop;
  reg _mul_6_source_busy;
  wire _mul_6_sink_start;
  wire _mul_6_sink_stop;
  wire _mul_6_sink_busy;
  wire _mul_6_busy;
  reg _mul_6_busy_reg;
  wire _mul_6_is_root;
  reg _mul_6_x_idle;
  reg [33-1:0] _mul_6_x_source_count;
  reg [5-1:0] _mul_6_x_source_mode;
  reg [16-1:0] _mul_6_x_source_generator_id;
  reg [32-1:0] _mul_6_x_source_offset;
  reg [33-1:0] _mul_6_x_source_size;
  reg [32-1:0] _mul_6_x_source_stride;
  reg [32-1:0] _mul_6_x_source_offset_buf;
  reg [33-1:0] _mul_6_x_source_size_buf;
  reg [32-1:0] _mul_6_x_source_stride_buf;
  reg [8-1:0] _mul_6_x_source_sel;
  reg [32-1:0] _mul_6_x_source_ram_raddr;
  reg _mul_6_x_source_ram_renable;
  wire [8-1:0] _mul_6_x_source_ram_rdata;
  reg _mul_6_x_source_fifo_deq;
  wire [8-1:0] _mul_6_x_source_fifo_rdata;
  reg [8-1:0] _mul_6_x_source_empty_data;
  reg _mul_6_y_idle;
  reg [33-1:0] _mul_6_y_source_count;
  reg [5-1:0] _mul_6_y_source_mode;
  reg [16-1:0] _mul_6_y_source_generator_id;
  reg [32-1:0] _mul_6_y_source_offset;
  reg [33-1:0] _mul_6_y_source_size;
  reg [32-1:0] _mul_6_y_source_stride;
  reg [32-1:0] _mul_6_y_source_offset_buf;
  reg [33-1:0] _mul_6_y_source_size_buf;
  reg [32-1:0] _mul_6_y_source_stride_buf;
  reg [8-1:0] _mul_6_y_source_sel;
  reg [32-1:0] _mul_6_y_source_ram_raddr;
  reg _mul_6_y_source_ram_renable;
  wire [8-1:0] _mul_6_y_source_ram_rdata;
  reg _mul_6_y_source_fifo_deq;
  wire [8-1:0] _mul_6_y_source_fifo_rdata;
  reg [8-1:0] _mul_6_y_source_empty_data;
  reg _mul_6_rshift_idle;
  reg [33-1:0] _mul_6_rshift_source_count;
  reg [5-1:0] _mul_6_rshift_source_mode;
  reg [16-1:0] _mul_6_rshift_source_generator_id;
  reg [32-1:0] _mul_6_rshift_source_offset;
  reg [33-1:0] _mul_6_rshift_source_size;
  reg [32-1:0] _mul_6_rshift_source_stride;
  reg [32-1:0] _mul_6_rshift_source_offset_buf;
  reg [33-1:0] _mul_6_rshift_source_size_buf;
  reg [32-1:0] _mul_6_rshift_source_stride_buf;
  reg [8-1:0] _mul_6_rshift_source_sel;
  reg [32-1:0] _mul_6_rshift_source_ram_raddr;
  reg _mul_6_rshift_source_ram_renable;
  wire [32-1:0] _mul_6_rshift_source_ram_rdata;
  reg _mul_6_rshift_source_fifo_deq;
  wire [32-1:0] _mul_6_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_6_rshift_source_empty_data;
  reg [33-1:0] _mul_6_z_sink_count;
  reg [5-1:0] _mul_6_z_sink_mode;
  reg [16-1:0] _mul_6_z_sink_generator_id;
  reg [32-1:0] _mul_6_z_sink_offset;
  reg [33-1:0] _mul_6_z_sink_size;
  reg [32-1:0] _mul_6_z_sink_stride;
  reg [32-1:0] _mul_6_z_sink_offset_buf;
  reg [33-1:0] _mul_6_z_sink_size_buf;
  reg [32-1:0] _mul_6_z_sink_stride_buf;
  reg [8-1:0] _mul_6_z_sink_sel;
  reg [32-1:0] _mul_6_z_sink_waddr;
  reg _mul_6_z_sink_wenable;
  reg [16-1:0] _mul_6_z_sink_wdata;
  reg _mul_6_z_sink_fifo_enq;
  reg [16-1:0] _mul_6_z_sink_fifo_wdata;
  reg [16-1:0] _mul_6_z_sink_immediate;
  reg _mul_7_stream_ivalid;
  wire _mul_7_stream_oready;
  wire _mul_7_stream_internal_oready;
  assign _mul_7_stream_internal_oready = 1;
  reg [32-1:0] _mul_7_fsm;
  localparam _mul_7_fsm_init = 0;
  wire _mul_7_run_flag;
  assign _mul_7_run_flag = 0;
  reg _mul_7_source_start;
  wire _mul_7_source_stop;
  reg _mul_7_source_busy;
  wire _mul_7_sink_start;
  wire _mul_7_sink_stop;
  wire _mul_7_sink_busy;
  wire _mul_7_busy;
  reg _mul_7_busy_reg;
  wire _mul_7_is_root;
  reg _mul_7_x_idle;
  reg [33-1:0] _mul_7_x_source_count;
  reg [5-1:0] _mul_7_x_source_mode;
  reg [16-1:0] _mul_7_x_source_generator_id;
  reg [32-1:0] _mul_7_x_source_offset;
  reg [33-1:0] _mul_7_x_source_size;
  reg [32-1:0] _mul_7_x_source_stride;
  reg [32-1:0] _mul_7_x_source_offset_buf;
  reg [33-1:0] _mul_7_x_source_size_buf;
  reg [32-1:0] _mul_7_x_source_stride_buf;
  reg [8-1:0] _mul_7_x_source_sel;
  reg [32-1:0] _mul_7_x_source_ram_raddr;
  reg _mul_7_x_source_ram_renable;
  wire [8-1:0] _mul_7_x_source_ram_rdata;
  reg _mul_7_x_source_fifo_deq;
  wire [8-1:0] _mul_7_x_source_fifo_rdata;
  reg [8-1:0] _mul_7_x_source_empty_data;
  reg _mul_7_y_idle;
  reg [33-1:0] _mul_7_y_source_count;
  reg [5-1:0] _mul_7_y_source_mode;
  reg [16-1:0] _mul_7_y_source_generator_id;
  reg [32-1:0] _mul_7_y_source_offset;
  reg [33-1:0] _mul_7_y_source_size;
  reg [32-1:0] _mul_7_y_source_stride;
  reg [32-1:0] _mul_7_y_source_offset_buf;
  reg [33-1:0] _mul_7_y_source_size_buf;
  reg [32-1:0] _mul_7_y_source_stride_buf;
  reg [8-1:0] _mul_7_y_source_sel;
  reg [32-1:0] _mul_7_y_source_ram_raddr;
  reg _mul_7_y_source_ram_renable;
  wire [8-1:0] _mul_7_y_source_ram_rdata;
  reg _mul_7_y_source_fifo_deq;
  wire [8-1:0] _mul_7_y_source_fifo_rdata;
  reg [8-1:0] _mul_7_y_source_empty_data;
  reg _mul_7_rshift_idle;
  reg [33-1:0] _mul_7_rshift_source_count;
  reg [5-1:0] _mul_7_rshift_source_mode;
  reg [16-1:0] _mul_7_rshift_source_generator_id;
  reg [32-1:0] _mul_7_rshift_source_offset;
  reg [33-1:0] _mul_7_rshift_source_size;
  reg [32-1:0] _mul_7_rshift_source_stride;
  reg [32-1:0] _mul_7_rshift_source_offset_buf;
  reg [33-1:0] _mul_7_rshift_source_size_buf;
  reg [32-1:0] _mul_7_rshift_source_stride_buf;
  reg [8-1:0] _mul_7_rshift_source_sel;
  reg [32-1:0] _mul_7_rshift_source_ram_raddr;
  reg _mul_7_rshift_source_ram_renable;
  wire [32-1:0] _mul_7_rshift_source_ram_rdata;
  reg _mul_7_rshift_source_fifo_deq;
  wire [32-1:0] _mul_7_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_7_rshift_source_empty_data;
  reg [33-1:0] _mul_7_z_sink_count;
  reg [5-1:0] _mul_7_z_sink_mode;
  reg [16-1:0] _mul_7_z_sink_generator_id;
  reg [32-1:0] _mul_7_z_sink_offset;
  reg [33-1:0] _mul_7_z_sink_size;
  reg [32-1:0] _mul_7_z_sink_stride;
  reg [32-1:0] _mul_7_z_sink_offset_buf;
  reg [33-1:0] _mul_7_z_sink_size_buf;
  reg [32-1:0] _mul_7_z_sink_stride_buf;
  reg [8-1:0] _mul_7_z_sink_sel;
  reg [32-1:0] _mul_7_z_sink_waddr;
  reg _mul_7_z_sink_wenable;
  reg [16-1:0] _mul_7_z_sink_wdata;
  reg _mul_7_z_sink_fifo_enq;
  reg [16-1:0] _mul_7_z_sink_fifo_wdata;
  reg [16-1:0] _mul_7_z_sink_immediate;
  reg _mul_8_stream_ivalid;
  wire _mul_8_stream_oready;
  wire _mul_8_stream_internal_oready;
  assign _mul_8_stream_internal_oready = 1;
  reg [32-1:0] _mul_8_fsm;
  localparam _mul_8_fsm_init = 0;
  wire _mul_8_run_flag;
  assign _mul_8_run_flag = 0;
  reg _mul_8_source_start;
  wire _mul_8_source_stop;
  reg _mul_8_source_busy;
  wire _mul_8_sink_start;
  wire _mul_8_sink_stop;
  wire _mul_8_sink_busy;
  wire _mul_8_busy;
  reg _mul_8_busy_reg;
  wire _mul_8_is_root;
  reg _mul_8_x_idle;
  reg [33-1:0] _mul_8_x_source_count;
  reg [5-1:0] _mul_8_x_source_mode;
  reg [16-1:0] _mul_8_x_source_generator_id;
  reg [32-1:0] _mul_8_x_source_offset;
  reg [33-1:0] _mul_8_x_source_size;
  reg [32-1:0] _mul_8_x_source_stride;
  reg [32-1:0] _mul_8_x_source_offset_buf;
  reg [33-1:0] _mul_8_x_source_size_buf;
  reg [32-1:0] _mul_8_x_source_stride_buf;
  reg [8-1:0] _mul_8_x_source_sel;
  reg [32-1:0] _mul_8_x_source_ram_raddr;
  reg _mul_8_x_source_ram_renable;
  wire [8-1:0] _mul_8_x_source_ram_rdata;
  reg _mul_8_x_source_fifo_deq;
  wire [8-1:0] _mul_8_x_source_fifo_rdata;
  reg [8-1:0] _mul_8_x_source_empty_data;
  reg _mul_8_y_idle;
  reg [33-1:0] _mul_8_y_source_count;
  reg [5-1:0] _mul_8_y_source_mode;
  reg [16-1:0] _mul_8_y_source_generator_id;
  reg [32-1:0] _mul_8_y_source_offset;
  reg [33-1:0] _mul_8_y_source_size;
  reg [32-1:0] _mul_8_y_source_stride;
  reg [32-1:0] _mul_8_y_source_offset_buf;
  reg [33-1:0] _mul_8_y_source_size_buf;
  reg [32-1:0] _mul_8_y_source_stride_buf;
  reg [8-1:0] _mul_8_y_source_sel;
  reg [32-1:0] _mul_8_y_source_ram_raddr;
  reg _mul_8_y_source_ram_renable;
  wire [8-1:0] _mul_8_y_source_ram_rdata;
  reg _mul_8_y_source_fifo_deq;
  wire [8-1:0] _mul_8_y_source_fifo_rdata;
  reg [8-1:0] _mul_8_y_source_empty_data;
  reg _mul_8_rshift_idle;
  reg [33-1:0] _mul_8_rshift_source_count;
  reg [5-1:0] _mul_8_rshift_source_mode;
  reg [16-1:0] _mul_8_rshift_source_generator_id;
  reg [32-1:0] _mul_8_rshift_source_offset;
  reg [33-1:0] _mul_8_rshift_source_size;
  reg [32-1:0] _mul_8_rshift_source_stride;
  reg [32-1:0] _mul_8_rshift_source_offset_buf;
  reg [33-1:0] _mul_8_rshift_source_size_buf;
  reg [32-1:0] _mul_8_rshift_source_stride_buf;
  reg [8-1:0] _mul_8_rshift_source_sel;
  reg [32-1:0] _mul_8_rshift_source_ram_raddr;
  reg _mul_8_rshift_source_ram_renable;
  wire [32-1:0] _mul_8_rshift_source_ram_rdata;
  reg _mul_8_rshift_source_fifo_deq;
  wire [32-1:0] _mul_8_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_8_rshift_source_empty_data;
  reg [33-1:0] _mul_8_z_sink_count;
  reg [5-1:0] _mul_8_z_sink_mode;
  reg [16-1:0] _mul_8_z_sink_generator_id;
  reg [32-1:0] _mul_8_z_sink_offset;
  reg [33-1:0] _mul_8_z_sink_size;
  reg [32-1:0] _mul_8_z_sink_stride;
  reg [32-1:0] _mul_8_z_sink_offset_buf;
  reg [33-1:0] _mul_8_z_sink_size_buf;
  reg [32-1:0] _mul_8_z_sink_stride_buf;
  reg [8-1:0] _mul_8_z_sink_sel;
  reg [32-1:0] _mul_8_z_sink_waddr;
  reg _mul_8_z_sink_wenable;
  reg [16-1:0] _mul_8_z_sink_wdata;
  reg _mul_8_z_sink_fifo_enq;
  reg [16-1:0] _mul_8_z_sink_fifo_wdata;
  reg [16-1:0] _mul_8_z_sink_immediate;
  reg _mul_9_stream_ivalid;
  wire _mul_9_stream_oready;
  wire _mul_9_stream_internal_oready;
  assign _mul_9_stream_internal_oready = 1;
  reg [32-1:0] _mul_9_fsm;
  localparam _mul_9_fsm_init = 0;
  wire _mul_9_run_flag;
  assign _mul_9_run_flag = 0;
  reg _mul_9_source_start;
  wire _mul_9_source_stop;
  reg _mul_9_source_busy;
  wire _mul_9_sink_start;
  wire _mul_9_sink_stop;
  wire _mul_9_sink_busy;
  wire _mul_9_busy;
  reg _mul_9_busy_reg;
  wire _mul_9_is_root;
  reg _mul_9_x_idle;
  reg [33-1:0] _mul_9_x_source_count;
  reg [5-1:0] _mul_9_x_source_mode;
  reg [16-1:0] _mul_9_x_source_generator_id;
  reg [32-1:0] _mul_9_x_source_offset;
  reg [33-1:0] _mul_9_x_source_size;
  reg [32-1:0] _mul_9_x_source_stride;
  reg [32-1:0] _mul_9_x_source_offset_buf;
  reg [33-1:0] _mul_9_x_source_size_buf;
  reg [32-1:0] _mul_9_x_source_stride_buf;
  reg [8-1:0] _mul_9_x_source_sel;
  reg [32-1:0] _mul_9_x_source_ram_raddr;
  reg _mul_9_x_source_ram_renable;
  wire [8-1:0] _mul_9_x_source_ram_rdata;
  reg _mul_9_x_source_fifo_deq;
  wire [8-1:0] _mul_9_x_source_fifo_rdata;
  reg [8-1:0] _mul_9_x_source_empty_data;
  reg _mul_9_y_idle;
  reg [33-1:0] _mul_9_y_source_count;
  reg [5-1:0] _mul_9_y_source_mode;
  reg [16-1:0] _mul_9_y_source_generator_id;
  reg [32-1:0] _mul_9_y_source_offset;
  reg [33-1:0] _mul_9_y_source_size;
  reg [32-1:0] _mul_9_y_source_stride;
  reg [32-1:0] _mul_9_y_source_offset_buf;
  reg [33-1:0] _mul_9_y_source_size_buf;
  reg [32-1:0] _mul_9_y_source_stride_buf;
  reg [8-1:0] _mul_9_y_source_sel;
  reg [32-1:0] _mul_9_y_source_ram_raddr;
  reg _mul_9_y_source_ram_renable;
  wire [8-1:0] _mul_9_y_source_ram_rdata;
  reg _mul_9_y_source_fifo_deq;
  wire [8-1:0] _mul_9_y_source_fifo_rdata;
  reg [8-1:0] _mul_9_y_source_empty_data;
  reg _mul_9_rshift_idle;
  reg [33-1:0] _mul_9_rshift_source_count;
  reg [5-1:0] _mul_9_rshift_source_mode;
  reg [16-1:0] _mul_9_rshift_source_generator_id;
  reg [32-1:0] _mul_9_rshift_source_offset;
  reg [33-1:0] _mul_9_rshift_source_size;
  reg [32-1:0] _mul_9_rshift_source_stride;
  reg [32-1:0] _mul_9_rshift_source_offset_buf;
  reg [33-1:0] _mul_9_rshift_source_size_buf;
  reg [32-1:0] _mul_9_rshift_source_stride_buf;
  reg [8-1:0] _mul_9_rshift_source_sel;
  reg [32-1:0] _mul_9_rshift_source_ram_raddr;
  reg _mul_9_rshift_source_ram_renable;
  wire [32-1:0] _mul_9_rshift_source_ram_rdata;
  reg _mul_9_rshift_source_fifo_deq;
  wire [32-1:0] _mul_9_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_9_rshift_source_empty_data;
  reg [33-1:0] _mul_9_z_sink_count;
  reg [5-1:0] _mul_9_z_sink_mode;
  reg [16-1:0] _mul_9_z_sink_generator_id;
  reg [32-1:0] _mul_9_z_sink_offset;
  reg [33-1:0] _mul_9_z_sink_size;
  reg [32-1:0] _mul_9_z_sink_stride;
  reg [32-1:0] _mul_9_z_sink_offset_buf;
  reg [33-1:0] _mul_9_z_sink_size_buf;
  reg [32-1:0] _mul_9_z_sink_stride_buf;
  reg [8-1:0] _mul_9_z_sink_sel;
  reg [32-1:0] _mul_9_z_sink_waddr;
  reg _mul_9_z_sink_wenable;
  reg [16-1:0] _mul_9_z_sink_wdata;
  reg _mul_9_z_sink_fifo_enq;
  reg [16-1:0] _mul_9_z_sink_fifo_wdata;
  reg [16-1:0] _mul_9_z_sink_immediate;
  reg _mul_10_stream_ivalid;
  wire _mul_10_stream_oready;
  wire _mul_10_stream_internal_oready;
  assign _mul_10_stream_internal_oready = 1;
  reg [32-1:0] _mul_10_fsm;
  localparam _mul_10_fsm_init = 0;
  wire _mul_10_run_flag;
  assign _mul_10_run_flag = 0;
  reg _mul_10_source_start;
  wire _mul_10_source_stop;
  reg _mul_10_source_busy;
  wire _mul_10_sink_start;
  wire _mul_10_sink_stop;
  wire _mul_10_sink_busy;
  wire _mul_10_busy;
  reg _mul_10_busy_reg;
  wire _mul_10_is_root;
  reg _mul_10_x_idle;
  reg [33-1:0] _mul_10_x_source_count;
  reg [5-1:0] _mul_10_x_source_mode;
  reg [16-1:0] _mul_10_x_source_generator_id;
  reg [32-1:0] _mul_10_x_source_offset;
  reg [33-1:0] _mul_10_x_source_size;
  reg [32-1:0] _mul_10_x_source_stride;
  reg [32-1:0] _mul_10_x_source_offset_buf;
  reg [33-1:0] _mul_10_x_source_size_buf;
  reg [32-1:0] _mul_10_x_source_stride_buf;
  reg [8-1:0] _mul_10_x_source_sel;
  reg [32-1:0] _mul_10_x_source_ram_raddr;
  reg _mul_10_x_source_ram_renable;
  wire [8-1:0] _mul_10_x_source_ram_rdata;
  reg _mul_10_x_source_fifo_deq;
  wire [8-1:0] _mul_10_x_source_fifo_rdata;
  reg [8-1:0] _mul_10_x_source_empty_data;
  reg _mul_10_y_idle;
  reg [33-1:0] _mul_10_y_source_count;
  reg [5-1:0] _mul_10_y_source_mode;
  reg [16-1:0] _mul_10_y_source_generator_id;
  reg [32-1:0] _mul_10_y_source_offset;
  reg [33-1:0] _mul_10_y_source_size;
  reg [32-1:0] _mul_10_y_source_stride;
  reg [32-1:0] _mul_10_y_source_offset_buf;
  reg [33-1:0] _mul_10_y_source_size_buf;
  reg [32-1:0] _mul_10_y_source_stride_buf;
  reg [8-1:0] _mul_10_y_source_sel;
  reg [32-1:0] _mul_10_y_source_ram_raddr;
  reg _mul_10_y_source_ram_renable;
  wire [8-1:0] _mul_10_y_source_ram_rdata;
  reg _mul_10_y_source_fifo_deq;
  wire [8-1:0] _mul_10_y_source_fifo_rdata;
  reg [8-1:0] _mul_10_y_source_empty_data;
  reg _mul_10_rshift_idle;
  reg [33-1:0] _mul_10_rshift_source_count;
  reg [5-1:0] _mul_10_rshift_source_mode;
  reg [16-1:0] _mul_10_rshift_source_generator_id;
  reg [32-1:0] _mul_10_rshift_source_offset;
  reg [33-1:0] _mul_10_rshift_source_size;
  reg [32-1:0] _mul_10_rshift_source_stride;
  reg [32-1:0] _mul_10_rshift_source_offset_buf;
  reg [33-1:0] _mul_10_rshift_source_size_buf;
  reg [32-1:0] _mul_10_rshift_source_stride_buf;
  reg [8-1:0] _mul_10_rshift_source_sel;
  reg [32-1:0] _mul_10_rshift_source_ram_raddr;
  reg _mul_10_rshift_source_ram_renable;
  wire [32-1:0] _mul_10_rshift_source_ram_rdata;
  reg _mul_10_rshift_source_fifo_deq;
  wire [32-1:0] _mul_10_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_10_rshift_source_empty_data;
  reg [33-1:0] _mul_10_z_sink_count;
  reg [5-1:0] _mul_10_z_sink_mode;
  reg [16-1:0] _mul_10_z_sink_generator_id;
  reg [32-1:0] _mul_10_z_sink_offset;
  reg [33-1:0] _mul_10_z_sink_size;
  reg [32-1:0] _mul_10_z_sink_stride;
  reg [32-1:0] _mul_10_z_sink_offset_buf;
  reg [33-1:0] _mul_10_z_sink_size_buf;
  reg [32-1:0] _mul_10_z_sink_stride_buf;
  reg [8-1:0] _mul_10_z_sink_sel;
  reg [32-1:0] _mul_10_z_sink_waddr;
  reg _mul_10_z_sink_wenable;
  reg [16-1:0] _mul_10_z_sink_wdata;
  reg _mul_10_z_sink_fifo_enq;
  reg [16-1:0] _mul_10_z_sink_fifo_wdata;
  reg [16-1:0] _mul_10_z_sink_immediate;
  reg _mul_11_stream_ivalid;
  wire _mul_11_stream_oready;
  wire _mul_11_stream_internal_oready;
  assign _mul_11_stream_internal_oready = 1;
  reg [32-1:0] _mul_11_fsm;
  localparam _mul_11_fsm_init = 0;
  wire _mul_11_run_flag;
  assign _mul_11_run_flag = 0;
  reg _mul_11_source_start;
  wire _mul_11_source_stop;
  reg _mul_11_source_busy;
  wire _mul_11_sink_start;
  wire _mul_11_sink_stop;
  wire _mul_11_sink_busy;
  wire _mul_11_busy;
  reg _mul_11_busy_reg;
  wire _mul_11_is_root;
  reg _mul_11_x_idle;
  reg [33-1:0] _mul_11_x_source_count;
  reg [5-1:0] _mul_11_x_source_mode;
  reg [16-1:0] _mul_11_x_source_generator_id;
  reg [32-1:0] _mul_11_x_source_offset;
  reg [33-1:0] _mul_11_x_source_size;
  reg [32-1:0] _mul_11_x_source_stride;
  reg [32-1:0] _mul_11_x_source_offset_buf;
  reg [33-1:0] _mul_11_x_source_size_buf;
  reg [32-1:0] _mul_11_x_source_stride_buf;
  reg [8-1:0] _mul_11_x_source_sel;
  reg [32-1:0] _mul_11_x_source_ram_raddr;
  reg _mul_11_x_source_ram_renable;
  wire [8-1:0] _mul_11_x_source_ram_rdata;
  reg _mul_11_x_source_fifo_deq;
  wire [8-1:0] _mul_11_x_source_fifo_rdata;
  reg [8-1:0] _mul_11_x_source_empty_data;
  reg _mul_11_y_idle;
  reg [33-1:0] _mul_11_y_source_count;
  reg [5-1:0] _mul_11_y_source_mode;
  reg [16-1:0] _mul_11_y_source_generator_id;
  reg [32-1:0] _mul_11_y_source_offset;
  reg [33-1:0] _mul_11_y_source_size;
  reg [32-1:0] _mul_11_y_source_stride;
  reg [32-1:0] _mul_11_y_source_offset_buf;
  reg [33-1:0] _mul_11_y_source_size_buf;
  reg [32-1:0] _mul_11_y_source_stride_buf;
  reg [8-1:0] _mul_11_y_source_sel;
  reg [32-1:0] _mul_11_y_source_ram_raddr;
  reg _mul_11_y_source_ram_renable;
  wire [8-1:0] _mul_11_y_source_ram_rdata;
  reg _mul_11_y_source_fifo_deq;
  wire [8-1:0] _mul_11_y_source_fifo_rdata;
  reg [8-1:0] _mul_11_y_source_empty_data;
  reg _mul_11_rshift_idle;
  reg [33-1:0] _mul_11_rshift_source_count;
  reg [5-1:0] _mul_11_rshift_source_mode;
  reg [16-1:0] _mul_11_rshift_source_generator_id;
  reg [32-1:0] _mul_11_rshift_source_offset;
  reg [33-1:0] _mul_11_rshift_source_size;
  reg [32-1:0] _mul_11_rshift_source_stride;
  reg [32-1:0] _mul_11_rshift_source_offset_buf;
  reg [33-1:0] _mul_11_rshift_source_size_buf;
  reg [32-1:0] _mul_11_rshift_source_stride_buf;
  reg [8-1:0] _mul_11_rshift_source_sel;
  reg [32-1:0] _mul_11_rshift_source_ram_raddr;
  reg _mul_11_rshift_source_ram_renable;
  wire [32-1:0] _mul_11_rshift_source_ram_rdata;
  reg _mul_11_rshift_source_fifo_deq;
  wire [32-1:0] _mul_11_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_11_rshift_source_empty_data;
  reg [33-1:0] _mul_11_z_sink_count;
  reg [5-1:0] _mul_11_z_sink_mode;
  reg [16-1:0] _mul_11_z_sink_generator_id;
  reg [32-1:0] _mul_11_z_sink_offset;
  reg [33-1:0] _mul_11_z_sink_size;
  reg [32-1:0] _mul_11_z_sink_stride;
  reg [32-1:0] _mul_11_z_sink_offset_buf;
  reg [33-1:0] _mul_11_z_sink_size_buf;
  reg [32-1:0] _mul_11_z_sink_stride_buf;
  reg [8-1:0] _mul_11_z_sink_sel;
  reg [32-1:0] _mul_11_z_sink_waddr;
  reg _mul_11_z_sink_wenable;
  reg [16-1:0] _mul_11_z_sink_wdata;
  reg _mul_11_z_sink_fifo_enq;
  reg [16-1:0] _mul_11_z_sink_fifo_wdata;
  reg [16-1:0] _mul_11_z_sink_immediate;
  reg _mul_12_stream_ivalid;
  wire _mul_12_stream_oready;
  wire _mul_12_stream_internal_oready;
  assign _mul_12_stream_internal_oready = 1;
  reg [32-1:0] _mul_12_fsm;
  localparam _mul_12_fsm_init = 0;
  wire _mul_12_run_flag;
  assign _mul_12_run_flag = 0;
  reg _mul_12_source_start;
  wire _mul_12_source_stop;
  reg _mul_12_source_busy;
  wire _mul_12_sink_start;
  wire _mul_12_sink_stop;
  wire _mul_12_sink_busy;
  wire _mul_12_busy;
  reg _mul_12_busy_reg;
  wire _mul_12_is_root;
  reg _mul_12_x_idle;
  reg [33-1:0] _mul_12_x_source_count;
  reg [5-1:0] _mul_12_x_source_mode;
  reg [16-1:0] _mul_12_x_source_generator_id;
  reg [32-1:0] _mul_12_x_source_offset;
  reg [33-1:0] _mul_12_x_source_size;
  reg [32-1:0] _mul_12_x_source_stride;
  reg [32-1:0] _mul_12_x_source_offset_buf;
  reg [33-1:0] _mul_12_x_source_size_buf;
  reg [32-1:0] _mul_12_x_source_stride_buf;
  reg [8-1:0] _mul_12_x_source_sel;
  reg [32-1:0] _mul_12_x_source_ram_raddr;
  reg _mul_12_x_source_ram_renable;
  wire [8-1:0] _mul_12_x_source_ram_rdata;
  reg _mul_12_x_source_fifo_deq;
  wire [8-1:0] _mul_12_x_source_fifo_rdata;
  reg [8-1:0] _mul_12_x_source_empty_data;
  reg _mul_12_y_idle;
  reg [33-1:0] _mul_12_y_source_count;
  reg [5-1:0] _mul_12_y_source_mode;
  reg [16-1:0] _mul_12_y_source_generator_id;
  reg [32-1:0] _mul_12_y_source_offset;
  reg [33-1:0] _mul_12_y_source_size;
  reg [32-1:0] _mul_12_y_source_stride;
  reg [32-1:0] _mul_12_y_source_offset_buf;
  reg [33-1:0] _mul_12_y_source_size_buf;
  reg [32-1:0] _mul_12_y_source_stride_buf;
  reg [8-1:0] _mul_12_y_source_sel;
  reg [32-1:0] _mul_12_y_source_ram_raddr;
  reg _mul_12_y_source_ram_renable;
  wire [8-1:0] _mul_12_y_source_ram_rdata;
  reg _mul_12_y_source_fifo_deq;
  wire [8-1:0] _mul_12_y_source_fifo_rdata;
  reg [8-1:0] _mul_12_y_source_empty_data;
  reg _mul_12_rshift_idle;
  reg [33-1:0] _mul_12_rshift_source_count;
  reg [5-1:0] _mul_12_rshift_source_mode;
  reg [16-1:0] _mul_12_rshift_source_generator_id;
  reg [32-1:0] _mul_12_rshift_source_offset;
  reg [33-1:0] _mul_12_rshift_source_size;
  reg [32-1:0] _mul_12_rshift_source_stride;
  reg [32-1:0] _mul_12_rshift_source_offset_buf;
  reg [33-1:0] _mul_12_rshift_source_size_buf;
  reg [32-1:0] _mul_12_rshift_source_stride_buf;
  reg [8-1:0] _mul_12_rshift_source_sel;
  reg [32-1:0] _mul_12_rshift_source_ram_raddr;
  reg _mul_12_rshift_source_ram_renable;
  wire [32-1:0] _mul_12_rshift_source_ram_rdata;
  reg _mul_12_rshift_source_fifo_deq;
  wire [32-1:0] _mul_12_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_12_rshift_source_empty_data;
  reg [33-1:0] _mul_12_z_sink_count;
  reg [5-1:0] _mul_12_z_sink_mode;
  reg [16-1:0] _mul_12_z_sink_generator_id;
  reg [32-1:0] _mul_12_z_sink_offset;
  reg [33-1:0] _mul_12_z_sink_size;
  reg [32-1:0] _mul_12_z_sink_stride;
  reg [32-1:0] _mul_12_z_sink_offset_buf;
  reg [33-1:0] _mul_12_z_sink_size_buf;
  reg [32-1:0] _mul_12_z_sink_stride_buf;
  reg [8-1:0] _mul_12_z_sink_sel;
  reg [32-1:0] _mul_12_z_sink_waddr;
  reg _mul_12_z_sink_wenable;
  reg [16-1:0] _mul_12_z_sink_wdata;
  reg _mul_12_z_sink_fifo_enq;
  reg [16-1:0] _mul_12_z_sink_fifo_wdata;
  reg [16-1:0] _mul_12_z_sink_immediate;
  reg _mul_13_stream_ivalid;
  wire _mul_13_stream_oready;
  wire _mul_13_stream_internal_oready;
  assign _mul_13_stream_internal_oready = 1;
  reg [32-1:0] _mul_13_fsm;
  localparam _mul_13_fsm_init = 0;
  wire _mul_13_run_flag;
  assign _mul_13_run_flag = 0;
  reg _mul_13_source_start;
  wire _mul_13_source_stop;
  reg _mul_13_source_busy;
  wire _mul_13_sink_start;
  wire _mul_13_sink_stop;
  wire _mul_13_sink_busy;
  wire _mul_13_busy;
  reg _mul_13_busy_reg;
  wire _mul_13_is_root;
  reg _mul_13_x_idle;
  reg [33-1:0] _mul_13_x_source_count;
  reg [5-1:0] _mul_13_x_source_mode;
  reg [16-1:0] _mul_13_x_source_generator_id;
  reg [32-1:0] _mul_13_x_source_offset;
  reg [33-1:0] _mul_13_x_source_size;
  reg [32-1:0] _mul_13_x_source_stride;
  reg [32-1:0] _mul_13_x_source_offset_buf;
  reg [33-1:0] _mul_13_x_source_size_buf;
  reg [32-1:0] _mul_13_x_source_stride_buf;
  reg [8-1:0] _mul_13_x_source_sel;
  reg [32-1:0] _mul_13_x_source_ram_raddr;
  reg _mul_13_x_source_ram_renable;
  wire [8-1:0] _mul_13_x_source_ram_rdata;
  reg _mul_13_x_source_fifo_deq;
  wire [8-1:0] _mul_13_x_source_fifo_rdata;
  reg [8-1:0] _mul_13_x_source_empty_data;
  reg _mul_13_y_idle;
  reg [33-1:0] _mul_13_y_source_count;
  reg [5-1:0] _mul_13_y_source_mode;
  reg [16-1:0] _mul_13_y_source_generator_id;
  reg [32-1:0] _mul_13_y_source_offset;
  reg [33-1:0] _mul_13_y_source_size;
  reg [32-1:0] _mul_13_y_source_stride;
  reg [32-1:0] _mul_13_y_source_offset_buf;
  reg [33-1:0] _mul_13_y_source_size_buf;
  reg [32-1:0] _mul_13_y_source_stride_buf;
  reg [8-1:0] _mul_13_y_source_sel;
  reg [32-1:0] _mul_13_y_source_ram_raddr;
  reg _mul_13_y_source_ram_renable;
  wire [8-1:0] _mul_13_y_source_ram_rdata;
  reg _mul_13_y_source_fifo_deq;
  wire [8-1:0] _mul_13_y_source_fifo_rdata;
  reg [8-1:0] _mul_13_y_source_empty_data;
  reg _mul_13_rshift_idle;
  reg [33-1:0] _mul_13_rshift_source_count;
  reg [5-1:0] _mul_13_rshift_source_mode;
  reg [16-1:0] _mul_13_rshift_source_generator_id;
  reg [32-1:0] _mul_13_rshift_source_offset;
  reg [33-1:0] _mul_13_rshift_source_size;
  reg [32-1:0] _mul_13_rshift_source_stride;
  reg [32-1:0] _mul_13_rshift_source_offset_buf;
  reg [33-1:0] _mul_13_rshift_source_size_buf;
  reg [32-1:0] _mul_13_rshift_source_stride_buf;
  reg [8-1:0] _mul_13_rshift_source_sel;
  reg [32-1:0] _mul_13_rshift_source_ram_raddr;
  reg _mul_13_rshift_source_ram_renable;
  wire [32-1:0] _mul_13_rshift_source_ram_rdata;
  reg _mul_13_rshift_source_fifo_deq;
  wire [32-1:0] _mul_13_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_13_rshift_source_empty_data;
  reg [33-1:0] _mul_13_z_sink_count;
  reg [5-1:0] _mul_13_z_sink_mode;
  reg [16-1:0] _mul_13_z_sink_generator_id;
  reg [32-1:0] _mul_13_z_sink_offset;
  reg [33-1:0] _mul_13_z_sink_size;
  reg [32-1:0] _mul_13_z_sink_stride;
  reg [32-1:0] _mul_13_z_sink_offset_buf;
  reg [33-1:0] _mul_13_z_sink_size_buf;
  reg [32-1:0] _mul_13_z_sink_stride_buf;
  reg [8-1:0] _mul_13_z_sink_sel;
  reg [32-1:0] _mul_13_z_sink_waddr;
  reg _mul_13_z_sink_wenable;
  reg [16-1:0] _mul_13_z_sink_wdata;
  reg _mul_13_z_sink_fifo_enq;
  reg [16-1:0] _mul_13_z_sink_fifo_wdata;
  reg [16-1:0] _mul_13_z_sink_immediate;
  reg __reduce_max_14_stream_ivalid;
  wire __reduce_max_14_stream_oready;
  wire __reduce_max_14_stream_internal_oready;
  assign __reduce_max_14_stream_internal_oready = 1;
  reg [32-1:0] __reduce_max_14_fsm;
  localparam __reduce_max_14_fsm_init = 0;
  wire __reduce_max_14_run_flag;
  assign __reduce_max_14_run_flag = 0;
  reg __reduce_max_14_source_start;
  wire __reduce_max_14_source_stop;
  reg __reduce_max_14_source_busy;
  wire __reduce_max_14_sink_start;
  wire __reduce_max_14_sink_stop;
  wire __reduce_max_14_sink_busy;
  wire __reduce_max_14_busy;
  reg __reduce_max_14_busy_reg;
  wire __reduce_max_14_is_root;
  reg __reduce_max_14_x_idle;
  reg [33-1:0] __reduce_max_14_x_source_count;
  reg [5-1:0] __reduce_max_14_x_source_mode;
  reg [16-1:0] __reduce_max_14_x_source_generator_id;
  reg [32-1:0] __reduce_max_14_x_source_offset;
  reg [33-1:0] __reduce_max_14_x_source_size;
  reg [32-1:0] __reduce_max_14_x_source_stride;
  reg [32-1:0] __reduce_max_14_x_source_offset_buf;
  reg [33-1:0] __reduce_max_14_x_source_size_buf;
  reg [32-1:0] __reduce_max_14_x_source_stride_buf;
  reg [8-1:0] __reduce_max_14_x_source_sel;
  reg [32-1:0] __reduce_max_14_x_source_ram_raddr;
  reg __reduce_max_14_x_source_ram_renable;
  wire [8-1:0] __reduce_max_14_x_source_ram_rdata;
  reg __reduce_max_14_x_source_fifo_deq;
  wire [8-1:0] __reduce_max_14_x_source_fifo_rdata;
  reg [8-1:0] __reduce_max_14_x_source_empty_data;
  reg [32-1:0] __reduce_max_14_size_next_parameter_data;
  reg [33-1:0] __reduce_max_14_data_sink_count;
  reg [5-1:0] __reduce_max_14_data_sink_mode;
  reg [16-1:0] __reduce_max_14_data_sink_generator_id;
  reg [32-1:0] __reduce_max_14_data_sink_offset;
  reg [33-1:0] __reduce_max_14_data_sink_size;
  reg [32-1:0] __reduce_max_14_data_sink_stride;
  reg [32-1:0] __reduce_max_14_data_sink_offset_buf;
  reg [33-1:0] __reduce_max_14_data_sink_size_buf;
  reg [32-1:0] __reduce_max_14_data_sink_stride_buf;
  reg [8-1:0] __reduce_max_14_data_sink_sel;
  reg [32-1:0] __reduce_max_14_data_sink_waddr;
  reg __reduce_max_14_data_sink_wenable;
  reg [8-1:0] __reduce_max_14_data_sink_wdata;
  reg __reduce_max_14_data_sink_fifo_enq;
  reg [8-1:0] __reduce_max_14_data_sink_fifo_wdata;
  reg [8-1:0] __reduce_max_14_data_sink_immediate;
  reg [33-1:0] __reduce_max_14_valid_sink_count;
  reg [5-1:0] __reduce_max_14_valid_sink_mode;
  reg [16-1:0] __reduce_max_14_valid_sink_generator_id;
  reg [32-1:0] __reduce_max_14_valid_sink_offset;
  reg [33-1:0] __reduce_max_14_valid_sink_size;
  reg [32-1:0] __reduce_max_14_valid_sink_stride;
  reg [32-1:0] __reduce_max_14_valid_sink_offset_buf;
  reg [33-1:0] __reduce_max_14_valid_sink_size_buf;
  reg [32-1:0] __reduce_max_14_valid_sink_stride_buf;
  reg [8-1:0] __reduce_max_14_valid_sink_sel;
  reg [32-1:0] __reduce_max_14_valid_sink_waddr;
  reg __reduce_max_14_valid_sink_wenable;
  reg [1-1:0] __reduce_max_14_valid_sink_wdata;
  reg __reduce_max_14_valid_sink_fifo_enq;
  reg [1-1:0] __reduce_max_14_valid_sink_fifo_wdata;
  reg [1-1:0] __reduce_max_14_valid_sink_immediate;
  reg _stream_conv2d_24_stream_ivalid;
  wire _stream_conv2d_24_stream_oready;
  wire _stream_conv2d_24_stream_internal_oready;
  assign _stream_conv2d_24_stream_oready = _stream_conv2d_24_stream_internal_oready;
  reg [32-1:0] _stream_conv2d_24_fsm;
  localparam _stream_conv2d_24_fsm_init = 0;
  wire _stream_conv2d_24_run_flag;
  reg _stream_conv2d_24_source_start;
  wire _stream_conv2d_24_source_stop;
  reg _stream_conv2d_24_source_busy;
  wire _stream_conv2d_24_sink_start;
  wire _stream_conv2d_24_sink_stop;
  wire _stream_conv2d_24_sink_busy;
  wire _stream_conv2d_24_busy;
  reg _stream_conv2d_24_busy_reg;
  wire _stream_conv2d_24_is_root;
  assign _stream_conv2d_24_is_root = 1;
  reg [10-1:0] _stream_conv2d_24_parameter_0_next_parameter_data;
  reg [2-1:0] _stream_conv2d_24_parameter_1_next_parameter_data;
  reg [2-1:0] _stream_conv2d_24_parameter_2_next_parameter_data;
  reg [9-1:0] _stream_conv2d_24_parameter_3_next_parameter_data;
  reg [1-1:0] _stream_conv2d_24_parameter_4_next_parameter_data;
  reg [1-1:0] _stream_conv2d_24_parameter_6_next_parameter_data;
  reg _stream_conv2d_24_source_7_idle;
  reg [33-1:0] _stream_conv2d_24_source_7_source_count;
  reg [5-1:0] _stream_conv2d_24_source_7_source_mode;
  reg [16-1:0] _stream_conv2d_24_source_7_source_generator_id;
  reg [32-1:0] _stream_conv2d_24_source_7_source_offset;
  reg [33-1:0] _stream_conv2d_24_source_7_source_size;
  reg [32-1:0] _stream_conv2d_24_source_7_source_stride;
  reg [32-1:0] _stream_conv2d_24_source_7_source_offset_buf;
  reg [33-1:0] _stream_conv2d_24_source_7_source_size_buf;
  reg [32-1:0] _stream_conv2d_24_source_7_source_stride_buf;
  reg [8-1:0] _stream_conv2d_24_source_7_source_sel;
  reg [32-1:0] _stream_conv2d_24_source_7_source_ram_raddr;
  reg _stream_conv2d_24_source_7_source_ram_renable;
  wire [32-1:0] _stream_conv2d_24_source_7_source_ram_rdata;
  reg _stream_conv2d_24_source_7_source_fifo_deq;
  wire [32-1:0] _stream_conv2d_24_source_7_source_fifo_rdata;
  reg [32-1:0] _stream_conv2d_24_source_7_source_empty_data;
  reg [1-1:0] _stream_conv2d_24_parameter_8_next_parameter_data;
  reg _stream_conv2d_24_source_9_idle;
  reg [33-1:0] _stream_conv2d_24_source_9_source_count;
  reg [5-1:0] _stream_conv2d_24_source_9_source_mode;
  reg [16-1:0] _stream_conv2d_24_source_9_source_generator_id;
  reg [32-1:0] _stream_conv2d_24_source_9_source_offset;
  reg [33-1:0] _stream_conv2d_24_source_9_source_size;
  reg [32-1:0] _stream_conv2d_24_source_9_source_stride;
  reg [32-1:0] _stream_conv2d_24_source_9_source_offset_buf;
  reg [33-1:0] _stream_conv2d_24_source_9_source_size_buf;
  reg [32-1:0] _stream_conv2d_24_source_9_source_stride_buf;
  reg [8-1:0] _stream_conv2d_24_source_9_source_sel;
  reg [32-1:0] _stream_conv2d_24_source_9_source_ram_raddr;
  reg _stream_conv2d_24_source_9_source_ram_renable;
  wire [8-1:0] _stream_conv2d_24_source_9_source_ram_rdata;
  reg _stream_conv2d_24_source_9_source_fifo_deq;
  wire [8-1:0] _stream_conv2d_24_source_9_source_fifo_rdata;
  reg [8-1:0] _stream_conv2d_24_source_9_source_empty_data;
  reg [1-1:0] _stream_conv2d_24_parameter_10_next_parameter_data;
  reg _stream_conv2d_24_source_11_idle;
  reg [33-1:0] _stream_conv2d_24_source_11_source_count;
  reg [5-1:0] _stream_conv2d_24_source_11_source_mode;
  reg [16-1:0] _stream_conv2d_24_source_11_source_generator_id;
  reg [32-1:0] _stream_conv2d_24_source_11_source_offset;
  reg [33-1:0] _stream_conv2d_24_source_11_source_size;
  reg [32-1:0] _stream_conv2d_24_source_11_source_stride;
  reg [32-1:0] _stream_conv2d_24_source_11_source_offset_buf;
  reg [33-1:0] _stream_conv2d_24_source_11_source_size_buf;
  reg [32-1:0] _stream_conv2d_24_source_11_source_stride_buf;
  reg [8-1:0] _stream_conv2d_24_source_11_source_sel;
  reg [32-1:0] _stream_conv2d_24_source_11_source_ram_raddr;
  reg _stream_conv2d_24_source_11_source_ram_renable;
  wire [8-1:0] _stream_conv2d_24_source_11_source_ram_rdata;
  reg _stream_conv2d_24_source_11_source_fifo_deq;
  wire [8-1:0] _stream_conv2d_24_source_11_source_fifo_rdata;
  reg [8-1:0] _stream_conv2d_24_source_11_source_empty_data;
  reg [1-1:0] _stream_conv2d_24_parameter_12_next_parameter_data;
  reg _stream_conv2d_24_source_13_idle;
  reg [33-1:0] _stream_conv2d_24_source_13_source_count;
  reg [5-1:0] _stream_conv2d_24_source_13_source_mode;
  reg [16-1:0] _stream_conv2d_24_source_13_source_generator_id;
  reg [32-1:0] _stream_conv2d_24_source_13_source_offset;
  reg [33-1:0] _stream_conv2d_24_source_13_source_size;
  reg [32-1:0] _stream_conv2d_24_source_13_source_stride;
  reg [32-1:0] _stream_conv2d_24_source_13_source_offset_buf;
  reg [33-1:0] _stream_conv2d_24_source_13_source_size_buf;
  reg [32-1:0] _stream_conv2d_24_source_13_source_stride_buf;
  reg [8-1:0] _stream_conv2d_24_source_13_source_sel;
  reg [32-1:0] _stream_conv2d_24_source_13_source_ram_raddr;
  reg _stream_conv2d_24_source_13_source_ram_renable;
  wire [8-1:0] _stream_conv2d_24_source_13_source_ram_rdata;
  reg _stream_conv2d_24_source_13_source_fifo_deq;
  wire [8-1:0] _stream_conv2d_24_source_13_source_fifo_rdata;
  reg [8-1:0] _stream_conv2d_24_source_13_source_empty_data;
  reg [1-1:0] _stream_conv2d_24_parameter_14_next_parameter_data;
  reg _stream_conv2d_24_source_15_idle;
  reg [33-1:0] _stream_conv2d_24_source_15_source_count;
  reg [5-1:0] _stream_conv2d_24_source_15_source_mode;
  reg [16-1:0] _stream_conv2d_24_source_15_source_generator_id;
  reg [32-1:0] _stream_conv2d_24_source_15_source_offset;
  reg [33-1:0] _stream_conv2d_24_source_15_source_size;
  reg [32-1:0] _stream_conv2d_24_source_15_source_stride;
  reg [32-1:0] _stream_conv2d_24_source_15_source_offset_buf;
  reg [33-1:0] _stream_conv2d_24_source_15_source_size_buf;
  reg [32-1:0] _stream_conv2d_24_source_15_source_stride_buf;
  reg [8-1:0] _stream_conv2d_24_source_15_source_sel;
  reg [32-1:0] _stream_conv2d_24_source_15_source_ram_raddr;
  reg _stream_conv2d_24_source_15_source_ram_renable;
  wire [8-1:0] _stream_conv2d_24_source_15_source_ram_rdata;
  reg _stream_conv2d_24_source_15_source_fifo_deq;
  wire [8-1:0] _stream_conv2d_24_source_15_source_fifo_rdata;
  reg [8-1:0] _stream_conv2d_24_source_15_source_empty_data;
  reg [1-1:0] _stream_conv2d_24_parameter_16_next_parameter_data;
  reg [1-1:0] _stream_conv2d_24_parameter_17_next_parameter_data;
  reg [5-1:0] _stream_conv2d_24_parameter_18_next_parameter_data;
  reg [1-1:0] _stream_conv2d_24_parameter_19_next_parameter_data;
  reg _stream_conv2d_24_source_20_idle;
  reg [33-1:0] _stream_conv2d_24_source_20_source_count;
  reg [5-1:0] _stream_conv2d_24_source_20_source_mode;
  reg [16-1:0] _stream_conv2d_24_source_20_source_generator_id;
  reg [32-1:0] _stream_conv2d_24_source_20_source_offset;
  reg [33-1:0] _stream_conv2d_24_source_20_source_size;
  reg [32-1:0] _stream_conv2d_24_source_20_source_stride;
  reg [32-1:0] _stream_conv2d_24_source_20_source_offset_buf;
  reg [33-1:0] _stream_conv2d_24_source_20_source_size_buf;
  reg [32-1:0] _stream_conv2d_24_source_20_source_stride_buf;
  reg [8-1:0] _stream_conv2d_24_source_20_source_sel;
  reg [32-1:0] _stream_conv2d_24_source_20_source_ram_raddr;
  reg _stream_conv2d_24_source_20_source_ram_renable;
  wire [8-1:0] _stream_conv2d_24_source_20_source_ram_rdata;
  reg _stream_conv2d_24_source_20_source_fifo_deq;
  wire [8-1:0] _stream_conv2d_24_source_20_source_fifo_rdata;
  reg [8-1:0] _stream_conv2d_24_source_20_source_empty_data;
  reg _stream_conv2d_24_source_21_idle;
  reg [33-1:0] _stream_conv2d_24_source_21_source_count;
  reg [5-1:0] _stream_conv2d_24_source_21_source_mode;
  reg [16-1:0] _stream_conv2d_24_source_21_source_generator_id;
  reg [32-1:0] _stream_conv2d_24_source_21_source_offset;
  reg [33-1:0] _stream_conv2d_24_source_21_source_size;
  reg [32-1:0] _stream_conv2d_24_source_21_source_stride;
  reg [32-1:0] _stream_conv2d_24_source_21_source_offset_buf;
  reg [33-1:0] _stream_conv2d_24_source_21_source_size_buf;
  reg [32-1:0] _stream_conv2d_24_source_21_source_stride_buf;
  reg [8-1:0] _stream_conv2d_24_source_21_source_sel;
  reg [32-1:0] _stream_conv2d_24_source_21_source_ram_raddr;
  reg _stream_conv2d_24_source_21_source_ram_renable;
  wire [8-1:0] _stream_conv2d_24_source_21_source_ram_rdata;
  reg _stream_conv2d_24_source_21_source_fifo_deq;
  wire [8-1:0] _stream_conv2d_24_source_21_source_fifo_rdata;
  reg [8-1:0] _stream_conv2d_24_source_21_source_empty_data;
  reg _stream_conv2d_24_source_22_idle;
  reg [33-1:0] _stream_conv2d_24_source_22_source_count;
  reg [5-1:0] _stream_conv2d_24_source_22_source_mode;
  reg [16-1:0] _stream_conv2d_24_source_22_source_generator_id;
  reg [32-1:0] _stream_conv2d_24_source_22_source_offset;
  reg [33-1:0] _stream_conv2d_24_source_22_source_size;
  reg [32-1:0] _stream_conv2d_24_source_22_source_stride;
  reg [32-1:0] _stream_conv2d_24_source_22_source_offset_buf;
  reg [33-1:0] _stream_conv2d_24_source_22_source_size_buf;
  reg [32-1:0] _stream_conv2d_24_source_22_source_stride_buf;
  reg [8-1:0] _stream_conv2d_24_source_22_source_sel;
  reg [32-1:0] _stream_conv2d_24_source_22_source_ram_raddr;
  reg _stream_conv2d_24_source_22_source_ram_renable;
  wire [8-1:0] _stream_conv2d_24_source_22_source_ram_rdata;
  reg _stream_conv2d_24_source_22_source_fifo_deq;
  wire [8-1:0] _stream_conv2d_24_source_22_source_fifo_rdata;
  reg [8-1:0] _stream_conv2d_24_source_22_source_empty_data;
  reg _stream_conv2d_24_source_23_idle;
  reg [33-1:0] _stream_conv2d_24_source_23_source_count;
  reg [5-1:0] _stream_conv2d_24_source_23_source_mode;
  reg [16-1:0] _stream_conv2d_24_source_23_source_generator_id;
  reg [32-1:0] _stream_conv2d_24_source_23_source_offset;
  reg [33-1:0] _stream_conv2d_24_source_23_source_size;
  reg [32-1:0] _stream_conv2d_24_source_23_source_stride;
  reg [32-1:0] _stream_conv2d_24_source_23_source_offset_buf;
  reg [33-1:0] _stream_conv2d_24_source_23_source_size_buf;
  reg [32-1:0] _stream_conv2d_24_source_23_source_stride_buf;
  reg [8-1:0] _stream_conv2d_24_source_23_source_sel;
  reg [32-1:0] _stream_conv2d_24_source_23_source_ram_raddr;
  reg _stream_conv2d_24_source_23_source_ram_renable;
  wire [8-1:0] _stream_conv2d_24_source_23_source_ram_rdata;
  reg _stream_conv2d_24_source_23_source_fifo_deq;
  wire [8-1:0] _stream_conv2d_24_source_23_source_fifo_rdata;
  reg [8-1:0] _stream_conv2d_24_source_23_source_empty_data;
  reg _stream_conv2d_24_source_24_idle;
  reg [33-1:0] _stream_conv2d_24_source_24_source_count;
  reg [5-1:0] _stream_conv2d_24_source_24_source_mode;
  reg [16-1:0] _stream_conv2d_24_source_24_source_generator_id;
  reg [32-1:0] _stream_conv2d_24_source_24_source_offset;
  reg [33-1:0] _stream_conv2d_24_source_24_source_size;
  reg [32-1:0] _stream_conv2d_24_source_24_source_stride;
  reg [32-1:0] _stream_conv2d_24_source_24_source_offset_buf;
  reg [33-1:0] _stream_conv2d_24_source_24_source_size_buf;
  reg [32-1:0] _stream_conv2d_24_source_24_source_stride_buf;
  reg [8-1:0] _stream_conv2d_24_source_24_source_sel;
  reg [32-1:0] _stream_conv2d_24_source_24_source_ram_raddr;
  reg _stream_conv2d_24_source_24_source_ram_renable;
  wire [8-1:0] _stream_conv2d_24_source_24_source_ram_rdata;
  reg _stream_conv2d_24_source_24_source_fifo_deq;
  wire [8-1:0] _stream_conv2d_24_source_24_source_fifo_rdata;
  reg [8-1:0] _stream_conv2d_24_source_24_source_empty_data;
  reg _stream_conv2d_24_source_25_idle;
  reg [33-1:0] _stream_conv2d_24_source_25_source_count;
  reg [5-1:0] _stream_conv2d_24_source_25_source_mode;
  reg [16-1:0] _stream_conv2d_24_source_25_source_generator_id;
  reg [32-1:0] _stream_conv2d_24_source_25_source_offset;
  reg [33-1:0] _stream_conv2d_24_source_25_source_size;
  reg [32-1:0] _stream_conv2d_24_source_25_source_stride;
  reg [32-1:0] _stream_conv2d_24_source_25_source_offset_buf;
  reg [33-1:0] _stream_conv2d_24_source_25_source_size_buf;
  reg [32-1:0] _stream_conv2d_24_source_25_source_stride_buf;
  reg [8-1:0] _stream_conv2d_24_source_25_source_sel;
  reg [32-1:0] _stream_conv2d_24_source_25_source_ram_raddr;
  reg _stream_conv2d_24_source_25_source_ram_renable;
  wire [8-1:0] _stream_conv2d_24_source_25_source_ram_rdata;
  reg _stream_conv2d_24_source_25_source_fifo_deq;
  wire [8-1:0] _stream_conv2d_24_source_25_source_fifo_rdata;
  reg [8-1:0] _stream_conv2d_24_source_25_source_empty_data;
  reg _stream_conv2d_24_source_26_idle;
  reg [33-1:0] _stream_conv2d_24_source_26_source_count;
  reg [5-1:0] _stream_conv2d_24_source_26_source_mode;
  reg [16-1:0] _stream_conv2d_24_source_26_source_generator_id;
  reg [32-1:0] _stream_conv2d_24_source_26_source_offset;
  reg [33-1:0] _stream_conv2d_24_source_26_source_size;
  reg [32-1:0] _stream_conv2d_24_source_26_source_stride;
  reg [32-1:0] _stream_conv2d_24_source_26_source_offset_buf;
  reg [33-1:0] _stream_conv2d_24_source_26_source_size_buf;
  reg [32-1:0] _stream_conv2d_24_source_26_source_stride_buf;
  reg [8-1:0] _stream_conv2d_24_source_26_source_sel;
  reg [32-1:0] _stream_conv2d_24_source_26_source_ram_raddr;
  reg _stream_conv2d_24_source_26_source_ram_renable;
  wire [8-1:0] _stream_conv2d_24_source_26_source_ram_rdata;
  reg _stream_conv2d_24_source_26_source_fifo_deq;
  wire [8-1:0] _stream_conv2d_24_source_26_source_fifo_rdata;
  reg [8-1:0] _stream_conv2d_24_source_26_source_empty_data;
  reg _stream_conv2d_24_source_27_idle;
  reg [33-1:0] _stream_conv2d_24_source_27_source_count;
  reg [5-1:0] _stream_conv2d_24_source_27_source_mode;
  reg [16-1:0] _stream_conv2d_24_source_27_source_generator_id;
  reg [32-1:0] _stream_conv2d_24_source_27_source_offset;
  reg [33-1:0] _stream_conv2d_24_source_27_source_size;
  reg [32-1:0] _stream_conv2d_24_source_27_source_stride;
  reg [32-1:0] _stream_conv2d_24_source_27_source_offset_buf;
  reg [33-1:0] _stream_conv2d_24_source_27_source_size_buf;
  reg [32-1:0] _stream_conv2d_24_source_27_source_stride_buf;
  reg [8-1:0] _stream_conv2d_24_source_27_source_sel;
  reg [32-1:0] _stream_conv2d_24_source_27_source_ram_raddr;
  reg _stream_conv2d_24_source_27_source_ram_renable;
  wire [8-1:0] _stream_conv2d_24_source_27_source_ram_rdata;
  reg _stream_conv2d_24_source_27_source_fifo_deq;
  wire [8-1:0] _stream_conv2d_24_source_27_source_fifo_rdata;
  reg [8-1:0] _stream_conv2d_24_source_27_source_empty_data;
  reg _stream_conv2d_24_source_28_idle;
  reg [33-1:0] _stream_conv2d_24_source_28_source_count;
  reg [5-1:0] _stream_conv2d_24_source_28_source_mode;
  reg [16-1:0] _stream_conv2d_24_source_28_source_generator_id;
  reg [32-1:0] _stream_conv2d_24_source_28_source_offset;
  reg [33-1:0] _stream_conv2d_24_source_28_source_size;
  reg [32-1:0] _stream_conv2d_24_source_28_source_stride;
  reg [32-1:0] _stream_conv2d_24_source_28_source_offset_buf;
  reg [33-1:0] _stream_conv2d_24_source_28_source_size_buf;
  reg [32-1:0] _stream_conv2d_24_source_28_source_stride_buf;
  reg [8-1:0] _stream_conv2d_24_source_28_source_sel;
  reg [32-1:0] _stream_conv2d_24_source_28_source_ram_raddr;
  reg _stream_conv2d_24_source_28_source_ram_renable;
  wire [8-1:0] _stream_conv2d_24_source_28_source_ram_rdata;
  reg _stream_conv2d_24_source_28_source_fifo_deq;
  wire [8-1:0] _stream_conv2d_24_source_28_source_fifo_rdata;
  reg [8-1:0] _stream_conv2d_24_source_28_source_empty_data;
  reg _stream_conv2d_24_source_29_idle;
  reg [33-1:0] _stream_conv2d_24_source_29_source_count;
  reg [5-1:0] _stream_conv2d_24_source_29_source_mode;
  reg [16-1:0] _stream_conv2d_24_source_29_source_generator_id;
  reg [32-1:0] _stream_conv2d_24_source_29_source_offset;
  reg [33-1:0] _stream_conv2d_24_source_29_source_size;
  reg [32-1:0] _stream_conv2d_24_source_29_source_stride;
  reg [32-1:0] _stream_conv2d_24_source_29_source_offset_buf;
  reg [33-1:0] _stream_conv2d_24_source_29_source_size_buf;
  reg [32-1:0] _stream_conv2d_24_source_29_source_stride_buf;
  reg [8-1:0] _stream_conv2d_24_source_29_source_sel;
  reg [32-1:0] _stream_conv2d_24_source_29_source_ram_raddr;
  reg _stream_conv2d_24_source_29_source_ram_renable;
  wire [8-1:0] _stream_conv2d_24_source_29_source_ram_rdata;
  reg _stream_conv2d_24_source_29_source_fifo_deq;
  wire [8-1:0] _stream_conv2d_24_source_29_source_fifo_rdata;
  reg [8-1:0] _stream_conv2d_24_source_29_source_empty_data;
  reg _stream_conv2d_24_source_30_idle;
  reg [33-1:0] _stream_conv2d_24_source_30_source_count;
  reg [5-1:0] _stream_conv2d_24_source_30_source_mode;
  reg [16-1:0] _stream_conv2d_24_source_30_source_generator_id;
  reg [32-1:0] _stream_conv2d_24_source_30_source_offset;
  reg [33-1:0] _stream_conv2d_24_source_30_source_size;
  reg [32-1:0] _stream_conv2d_24_source_30_source_stride;
  reg [32-1:0] _stream_conv2d_24_source_30_source_offset_buf;
  reg [33-1:0] _stream_conv2d_24_source_30_source_size_buf;
  reg [32-1:0] _stream_conv2d_24_source_30_source_stride_buf;
  reg [8-1:0] _stream_conv2d_24_source_30_source_sel;
  reg [32-1:0] _stream_conv2d_24_source_30_source_ram_raddr;
  reg _stream_conv2d_24_source_30_source_ram_renable;
  wire [8-1:0] _stream_conv2d_24_source_30_source_ram_rdata;
  reg _stream_conv2d_24_source_30_source_fifo_deq;
  wire [8-1:0] _stream_conv2d_24_source_30_source_fifo_rdata;
  reg [8-1:0] _stream_conv2d_24_source_30_source_empty_data;
  reg _stream_conv2d_24_source_31_idle;
  reg [33-1:0] _stream_conv2d_24_source_31_source_count;
  reg [5-1:0] _stream_conv2d_24_source_31_source_mode;
  reg [16-1:0] _stream_conv2d_24_source_31_source_generator_id;
  reg [32-1:0] _stream_conv2d_24_source_31_source_offset;
  reg [33-1:0] _stream_conv2d_24_source_31_source_size;
  reg [32-1:0] _stream_conv2d_24_source_31_source_stride;
  reg [32-1:0] _stream_conv2d_24_source_31_source_offset_buf;
  reg [33-1:0] _stream_conv2d_24_source_31_source_size_buf;
  reg [32-1:0] _stream_conv2d_24_source_31_source_stride_buf;
  reg [8-1:0] _stream_conv2d_24_source_31_source_sel;
  reg [32-1:0] _stream_conv2d_24_source_31_source_ram_raddr;
  reg _stream_conv2d_24_source_31_source_ram_renable;
  wire [8-1:0] _stream_conv2d_24_source_31_source_ram_rdata;
  reg _stream_conv2d_24_source_31_source_fifo_deq;
  wire [8-1:0] _stream_conv2d_24_source_31_source_fifo_rdata;
  reg [8-1:0] _stream_conv2d_24_source_31_source_empty_data;
  reg _stream_conv2d_24_source_32_idle;
  reg [33-1:0] _stream_conv2d_24_source_32_source_count;
  reg [5-1:0] _stream_conv2d_24_source_32_source_mode;
  reg [16-1:0] _stream_conv2d_24_source_32_source_generator_id;
  reg [32-1:0] _stream_conv2d_24_source_32_source_offset;
  reg [33-1:0] _stream_conv2d_24_source_32_source_size;
  reg [32-1:0] _stream_conv2d_24_source_32_source_stride;
  reg [32-1:0] _stream_conv2d_24_source_32_source_offset_buf;
  reg [33-1:0] _stream_conv2d_24_source_32_source_size_buf;
  reg [32-1:0] _stream_conv2d_24_source_32_source_stride_buf;
  reg [8-1:0] _stream_conv2d_24_source_32_source_sel;
  reg [32-1:0] _stream_conv2d_24_source_32_source_ram_raddr;
  reg _stream_conv2d_24_source_32_source_ram_renable;
  wire [8-1:0] _stream_conv2d_24_source_32_source_ram_rdata;
  reg _stream_conv2d_24_source_32_source_fifo_deq;
  wire [8-1:0] _stream_conv2d_24_source_32_source_fifo_rdata;
  reg [8-1:0] _stream_conv2d_24_source_32_source_empty_data;
  reg _stream_conv2d_24_source_33_idle;
  reg [33-1:0] _stream_conv2d_24_source_33_source_count;
  reg [5-1:0] _stream_conv2d_24_source_33_source_mode;
  reg [16-1:0] _stream_conv2d_24_source_33_source_generator_id;
  reg [32-1:0] _stream_conv2d_24_source_33_source_offset;
  reg [33-1:0] _stream_conv2d_24_source_33_source_size;
  reg [32-1:0] _stream_conv2d_24_source_33_source_stride;
  reg [32-1:0] _stream_conv2d_24_source_33_source_offset_buf;
  reg [33-1:0] _stream_conv2d_24_source_33_source_size_buf;
  reg [32-1:0] _stream_conv2d_24_source_33_source_stride_buf;
  reg [8-1:0] _stream_conv2d_24_source_33_source_sel;
  reg [32-1:0] _stream_conv2d_24_source_33_source_ram_raddr;
  reg _stream_conv2d_24_source_33_source_ram_renable;
  wire [8-1:0] _stream_conv2d_24_source_33_source_ram_rdata;
  reg _stream_conv2d_24_source_33_source_fifo_deq;
  wire [8-1:0] _stream_conv2d_24_source_33_source_fifo_rdata;
  reg [8-1:0] _stream_conv2d_24_source_33_source_empty_data;
  reg _stream_conv2d_24_source_34_idle;
  reg [33-1:0] _stream_conv2d_24_source_34_source_count;
  reg [5-1:0] _stream_conv2d_24_source_34_source_mode;
  reg [16-1:0] _stream_conv2d_24_source_34_source_generator_id;
  reg [32-1:0] _stream_conv2d_24_source_34_source_offset;
  reg [33-1:0] _stream_conv2d_24_source_34_source_size;
  reg [32-1:0] _stream_conv2d_24_source_34_source_stride;
  reg [32-1:0] _stream_conv2d_24_source_34_source_offset_buf;
  reg [33-1:0] _stream_conv2d_24_source_34_source_size_buf;
  reg [32-1:0] _stream_conv2d_24_source_34_source_stride_buf;
  reg [8-1:0] _stream_conv2d_24_source_34_source_sel;
  reg [32-1:0] _stream_conv2d_24_source_34_source_ram_raddr;
  reg _stream_conv2d_24_source_34_source_ram_renable;
  wire [8-1:0] _stream_conv2d_24_source_34_source_ram_rdata;
  reg _stream_conv2d_24_source_34_source_fifo_deq;
  wire [8-1:0] _stream_conv2d_24_source_34_source_fifo_rdata;
  reg [8-1:0] _stream_conv2d_24_source_34_source_empty_data;
  reg _stream_conv2d_24_source_35_idle;
  reg [33-1:0] _stream_conv2d_24_source_35_source_count;
  reg [5-1:0] _stream_conv2d_24_source_35_source_mode;
  reg [16-1:0] _stream_conv2d_24_source_35_source_generator_id;
  reg [32-1:0] _stream_conv2d_24_source_35_source_offset;
  reg [33-1:0] _stream_conv2d_24_source_35_source_size;
  reg [32-1:0] _stream_conv2d_24_source_35_source_stride;
  reg [32-1:0] _stream_conv2d_24_source_35_source_offset_buf;
  reg [33-1:0] _stream_conv2d_24_source_35_source_size_buf;
  reg [32-1:0] _stream_conv2d_24_source_35_source_stride_buf;
  reg [8-1:0] _stream_conv2d_24_source_35_source_sel;
  reg [32-1:0] _stream_conv2d_24_source_35_source_ram_raddr;
  reg _stream_conv2d_24_source_35_source_ram_renable;
  wire [8-1:0] _stream_conv2d_24_source_35_source_ram_rdata;
  reg _stream_conv2d_24_source_35_source_fifo_deq;
  wire [8-1:0] _stream_conv2d_24_source_35_source_fifo_rdata;
  reg [8-1:0] _stream_conv2d_24_source_35_source_empty_data;
  reg _stream_conv2d_24_source_36_idle;
  reg [33-1:0] _stream_conv2d_24_source_36_source_count;
  reg [5-1:0] _stream_conv2d_24_source_36_source_mode;
  reg [16-1:0] _stream_conv2d_24_source_36_source_generator_id;
  reg [32-1:0] _stream_conv2d_24_source_36_source_offset;
  reg [33-1:0] _stream_conv2d_24_source_36_source_size;
  reg [32-1:0] _stream_conv2d_24_source_36_source_stride;
  reg [32-1:0] _stream_conv2d_24_source_36_source_offset_buf;
  reg [33-1:0] _stream_conv2d_24_source_36_source_size_buf;
  reg [32-1:0] _stream_conv2d_24_source_36_source_stride_buf;
  reg [8-1:0] _stream_conv2d_24_source_36_source_sel;
  reg [32-1:0] _stream_conv2d_24_source_36_source_ram_raddr;
  reg _stream_conv2d_24_source_36_source_ram_renable;
  wire [8-1:0] _stream_conv2d_24_source_36_source_ram_rdata;
  reg _stream_conv2d_24_source_36_source_fifo_deq;
  wire [8-1:0] _stream_conv2d_24_source_36_source_fifo_rdata;
  reg [8-1:0] _stream_conv2d_24_source_36_source_empty_data;
  reg _stream_conv2d_24_source_37_idle;
  reg [33-1:0] _stream_conv2d_24_source_37_source_count;
  reg [5-1:0] _stream_conv2d_24_source_37_source_mode;
  reg [16-1:0] _stream_conv2d_24_source_37_source_generator_id;
  reg [32-1:0] _stream_conv2d_24_source_37_source_offset;
  reg [33-1:0] _stream_conv2d_24_source_37_source_size;
  reg [32-1:0] _stream_conv2d_24_source_37_source_stride;
  reg [32-1:0] _stream_conv2d_24_source_37_source_offset_buf;
  reg [33-1:0] _stream_conv2d_24_source_37_source_size_buf;
  reg [32-1:0] _stream_conv2d_24_source_37_source_stride_buf;
  reg [8-1:0] _stream_conv2d_24_source_37_source_sel;
  reg [32-1:0] _stream_conv2d_24_source_37_source_ram_raddr;
  reg _stream_conv2d_24_source_37_source_ram_renable;
  wire [8-1:0] _stream_conv2d_24_source_37_source_ram_rdata;
  reg _stream_conv2d_24_source_37_source_fifo_deq;
  wire [8-1:0] _stream_conv2d_24_source_37_source_fifo_rdata;
  reg [8-1:0] _stream_conv2d_24_source_37_source_empty_data;
  wire signed [8-1:0] mul_5_x_data;
  wire signed [8-1:0] mul_5_y_data;
  wire [4-1:0] mul_5_rshift_data;
  reg __mul_5_stream_ivalid_1;
  reg __mul_5_stream_ivalid_2;
  reg __mul_5_stream_ivalid_3;
  reg __mul_5_stream_ivalid_4;
  reg __mul_5_stream_ivalid_5;
  reg __mul_5_stream_ivalid_6;
  reg __mul_5_stream_ivalid_7;
  reg __mul_5_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_111;
  reg [4-1:0] _minus_data_113;
  reg [1-1:0] _greatereq_data_124;
  reg signed [8-1:0] __delay_data_686__variable_108;
  reg signed [8-1:0] __delay_data_689__variable_109;
  reg [4-1:0] __delay_data_692__variable_110;
  reg signed [18-1:0] _sll_data_115;
  reg [1-1:0] __delay_data_683_greaterthan_111;
  reg [1-1:0] __delay_data_684_greatereq_124;
  reg signed [8-1:0] __delay_data_687__delay_686__variable_108;
  reg signed [8-1:0] __delay_data_690__delay_689__variable_109;
  reg [4-1:0] __delay_data_693__delay_692__variable_110;
  reg signed [16-1:0] _cond_data_121;
  reg [1-1:0] __delay_data_685__delay_684_greatereq_124;
  reg signed [8-1:0] __delay_data_688__delay_687__delay_686__variable_108;
  reg signed [8-1:0] __delay_data_691__delay_690__delay_689__variable_109;
  reg [4-1:0] __delay_data_694__delay_693__delay_692__variable_110;
  wire signed [8-1:0] _uminus_data_123;
  assign _uminus_data_123 = -_cond_data_121;
  wire signed [8-1:0] _cond_data_126;
  assign _cond_data_126 = (__delay_data_685__delay_684_greatereq_124)? _cond_data_121 : _uminus_data_123;
  wire signed [16-1:0] __muladd_madd_odata_127;
  reg signed [16-1:0] __muladd_madd_odata_reg_127;
  wire signed [16-1:0] __muladd_data_127;
  assign __muladd_data_127 = __muladd_madd_odata_reg_127;
  wire __muladd_madd_update_127;
  assign __muladd_madd_update_127 = _mul_5_stream_oready;

  madd_0
  __muladd_madd_127
  (
    .CLK(CLK),
    .update(__muladd_madd_update_127),
    .a(__delay_data_688__delay_687__delay_686__variable_108),
    .b(__delay_data_691__delay_690__delay_689__variable_109),
    .c(_cond_data_126),
    .d(__muladd_madd_odata_127)
  );

  reg [4-1:0] __delay_data_695__delay_694__delay_693____variable_110;
  reg [4-1:0] __delay_data_696__delay_695__delay_694____variable_110;
  reg [4-1:0] __delay_data_697__delay_696__delay_695____variable_110;
  reg [4-1:0] __delay_data_698__delay_697__delay_696____variable_110;
  reg signed [16-1:0] _sra_data_128;
  wire signed [16-1:0] mul_5_z_data;
  assign mul_5_z_data = _sra_data_128;
  wire signed [8-1:0] mul_6_x_data;
  wire signed [8-1:0] mul_6_y_data;
  wire [4-1:0] mul_6_rshift_data;
  reg __mul_6_stream_ivalid_1;
  reg __mul_6_stream_ivalid_2;
  reg __mul_6_stream_ivalid_3;
  reg __mul_6_stream_ivalid_4;
  reg __mul_6_stream_ivalid_5;
  reg __mul_6_stream_ivalid_6;
  reg __mul_6_stream_ivalid_7;
  reg __mul_6_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_132;
  reg [4-1:0] _minus_data_134;
  reg [1-1:0] _greatereq_data_145;
  reg signed [8-1:0] __delay_data_705__variable_129;
  reg signed [8-1:0] __delay_data_708__variable_130;
  reg [4-1:0] __delay_data_711__variable_131;
  reg signed [18-1:0] _sll_data_136;
  reg [1-1:0] __delay_data_702_greaterthan_132;
  reg [1-1:0] __delay_data_703_greatereq_145;
  reg signed [8-1:0] __delay_data_706__delay_705__variable_129;
  reg signed [8-1:0] __delay_data_709__delay_708__variable_130;
  reg [4-1:0] __delay_data_712__delay_711__variable_131;
  reg signed [16-1:0] _cond_data_142;
  reg [1-1:0] __delay_data_704__delay_703_greatereq_145;
  reg signed [8-1:0] __delay_data_707__delay_706__delay_705__variable_129;
  reg signed [8-1:0] __delay_data_710__delay_709__delay_708__variable_130;
  reg [4-1:0] __delay_data_713__delay_712__delay_711__variable_131;
  wire signed [8-1:0] _uminus_data_144;
  assign _uminus_data_144 = -_cond_data_142;
  wire signed [8-1:0] _cond_data_147;
  assign _cond_data_147 = (__delay_data_704__delay_703_greatereq_145)? _cond_data_142 : _uminus_data_144;
  wire signed [16-1:0] __muladd_madd_odata_148;
  reg signed [16-1:0] __muladd_madd_odata_reg_148;
  wire signed [16-1:0] __muladd_data_148;
  assign __muladd_data_148 = __muladd_madd_odata_reg_148;
  wire __muladd_madd_update_148;
  assign __muladd_madd_update_148 = _mul_6_stream_oready;

  madd_1
  __muladd_madd_148
  (
    .CLK(CLK),
    .update(__muladd_madd_update_148),
    .a(__delay_data_707__delay_706__delay_705__variable_129),
    .b(__delay_data_710__delay_709__delay_708__variable_130),
    .c(_cond_data_147),
    .d(__muladd_madd_odata_148)
  );

  reg [4-1:0] __delay_data_714__delay_713__delay_712____variable_131;
  reg [4-1:0] __delay_data_715__delay_714__delay_713____variable_131;
  reg [4-1:0] __delay_data_716__delay_715__delay_714____variable_131;
  reg [4-1:0] __delay_data_717__delay_716__delay_715____variable_131;
  reg signed [16-1:0] _sra_data_149;
  wire signed [16-1:0] mul_6_z_data;
  assign mul_6_z_data = _sra_data_149;
  wire signed [8-1:0] mul_7_x_data;
  wire signed [8-1:0] mul_7_y_data;
  wire [4-1:0] mul_7_rshift_data;
  reg __mul_7_stream_ivalid_1;
  reg __mul_7_stream_ivalid_2;
  reg __mul_7_stream_ivalid_3;
  reg __mul_7_stream_ivalid_4;
  reg __mul_7_stream_ivalid_5;
  reg __mul_7_stream_ivalid_6;
  reg __mul_7_stream_ivalid_7;
  reg __mul_7_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_153;
  reg [4-1:0] _minus_data_155;
  reg [1-1:0] _greatereq_data_166;
  reg signed [8-1:0] __delay_data_724__variable_150;
  reg signed [8-1:0] __delay_data_727__variable_151;
  reg [4-1:0] __delay_data_730__variable_152;
  reg signed [18-1:0] _sll_data_157;
  reg [1-1:0] __delay_data_721_greaterthan_153;
  reg [1-1:0] __delay_data_722_greatereq_166;
  reg signed [8-1:0] __delay_data_725__delay_724__variable_150;
  reg signed [8-1:0] __delay_data_728__delay_727__variable_151;
  reg [4-1:0] __delay_data_731__delay_730__variable_152;
  reg signed [16-1:0] _cond_data_163;
  reg [1-1:0] __delay_data_723__delay_722_greatereq_166;
  reg signed [8-1:0] __delay_data_726__delay_725__delay_724__variable_150;
  reg signed [8-1:0] __delay_data_729__delay_728__delay_727__variable_151;
  reg [4-1:0] __delay_data_732__delay_731__delay_730__variable_152;
  wire signed [8-1:0] _uminus_data_165;
  assign _uminus_data_165 = -_cond_data_163;
  wire signed [8-1:0] _cond_data_168;
  assign _cond_data_168 = (__delay_data_723__delay_722_greatereq_166)? _cond_data_163 : _uminus_data_165;
  wire signed [16-1:0] __muladd_madd_odata_169;
  reg signed [16-1:0] __muladd_madd_odata_reg_169;
  wire signed [16-1:0] __muladd_data_169;
  assign __muladd_data_169 = __muladd_madd_odata_reg_169;
  wire __muladd_madd_update_169;
  assign __muladd_madd_update_169 = _mul_7_stream_oready;

  madd_2
  __muladd_madd_169
  (
    .CLK(CLK),
    .update(__muladd_madd_update_169),
    .a(__delay_data_726__delay_725__delay_724__variable_150),
    .b(__delay_data_729__delay_728__delay_727__variable_151),
    .c(_cond_data_168),
    .d(__muladd_madd_odata_169)
  );

  reg [4-1:0] __delay_data_733__delay_732__delay_731____variable_152;
  reg [4-1:0] __delay_data_734__delay_733__delay_732____variable_152;
  reg [4-1:0] __delay_data_735__delay_734__delay_733____variable_152;
  reg [4-1:0] __delay_data_736__delay_735__delay_734____variable_152;
  reg signed [16-1:0] _sra_data_170;
  wire signed [16-1:0] mul_7_z_data;
  assign mul_7_z_data = _sra_data_170;
  wire signed [8-1:0] mul_8_x_data;
  wire signed [8-1:0] mul_8_y_data;
  wire [4-1:0] mul_8_rshift_data;
  reg __mul_8_stream_ivalid_1;
  reg __mul_8_stream_ivalid_2;
  reg __mul_8_stream_ivalid_3;
  reg __mul_8_stream_ivalid_4;
  reg __mul_8_stream_ivalid_5;
  reg __mul_8_stream_ivalid_6;
  reg __mul_8_stream_ivalid_7;
  reg __mul_8_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_174;
  reg [4-1:0] _minus_data_176;
  reg [1-1:0] _greatereq_data_187;
  reg signed [8-1:0] __delay_data_743__variable_171;
  reg signed [8-1:0] __delay_data_746__variable_172;
  reg [4-1:0] __delay_data_749__variable_173;
  reg signed [18-1:0] _sll_data_178;
  reg [1-1:0] __delay_data_740_greaterthan_174;
  reg [1-1:0] __delay_data_741_greatereq_187;
  reg signed [8-1:0] __delay_data_744__delay_743__variable_171;
  reg signed [8-1:0] __delay_data_747__delay_746__variable_172;
  reg [4-1:0] __delay_data_750__delay_749__variable_173;
  reg signed [16-1:0] _cond_data_184;
  reg [1-1:0] __delay_data_742__delay_741_greatereq_187;
  reg signed [8-1:0] __delay_data_745__delay_744__delay_743__variable_171;
  reg signed [8-1:0] __delay_data_748__delay_747__delay_746__variable_172;
  reg [4-1:0] __delay_data_751__delay_750__delay_749__variable_173;
  wire signed [8-1:0] _uminus_data_186;
  assign _uminus_data_186 = -_cond_data_184;
  wire signed [8-1:0] _cond_data_189;
  assign _cond_data_189 = (__delay_data_742__delay_741_greatereq_187)? _cond_data_184 : _uminus_data_186;
  wire signed [16-1:0] __muladd_madd_odata_190;
  reg signed [16-1:0] __muladd_madd_odata_reg_190;
  wire signed [16-1:0] __muladd_data_190;
  assign __muladd_data_190 = __muladd_madd_odata_reg_190;
  wire __muladd_madd_update_190;
  assign __muladd_madd_update_190 = _mul_8_stream_oready;

  madd_3
  __muladd_madd_190
  (
    .CLK(CLK),
    .update(__muladd_madd_update_190),
    .a(__delay_data_745__delay_744__delay_743__variable_171),
    .b(__delay_data_748__delay_747__delay_746__variable_172),
    .c(_cond_data_189),
    .d(__muladd_madd_odata_190)
  );

  reg [4-1:0] __delay_data_752__delay_751__delay_750____variable_173;
  reg [4-1:0] __delay_data_753__delay_752__delay_751____variable_173;
  reg [4-1:0] __delay_data_754__delay_753__delay_752____variable_173;
  reg [4-1:0] __delay_data_755__delay_754__delay_753____variable_173;
  reg signed [16-1:0] _sra_data_191;
  wire signed [16-1:0] mul_8_z_data;
  assign mul_8_z_data = _sra_data_191;
  wire signed [8-1:0] mul_9_x_data;
  wire signed [8-1:0] mul_9_y_data;
  wire [4-1:0] mul_9_rshift_data;
  reg __mul_9_stream_ivalid_1;
  reg __mul_9_stream_ivalid_2;
  reg __mul_9_stream_ivalid_3;
  reg __mul_9_stream_ivalid_4;
  reg __mul_9_stream_ivalid_5;
  reg __mul_9_stream_ivalid_6;
  reg __mul_9_stream_ivalid_7;
  reg __mul_9_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_195;
  reg [4-1:0] _minus_data_197;
  reg [1-1:0] _greatereq_data_208;
  reg signed [8-1:0] __delay_data_762__variable_192;
  reg signed [8-1:0] __delay_data_765__variable_193;
  reg [4-1:0] __delay_data_768__variable_194;
  reg signed [18-1:0] _sll_data_199;
  reg [1-1:0] __delay_data_759_greaterthan_195;
  reg [1-1:0] __delay_data_760_greatereq_208;
  reg signed [8-1:0] __delay_data_763__delay_762__variable_192;
  reg signed [8-1:0] __delay_data_766__delay_765__variable_193;
  reg [4-1:0] __delay_data_769__delay_768__variable_194;
  reg signed [16-1:0] _cond_data_205;
  reg [1-1:0] __delay_data_761__delay_760_greatereq_208;
  reg signed [8-1:0] __delay_data_764__delay_763__delay_762__variable_192;
  reg signed [8-1:0] __delay_data_767__delay_766__delay_765__variable_193;
  reg [4-1:0] __delay_data_770__delay_769__delay_768__variable_194;
  wire signed [8-1:0] _uminus_data_207;
  assign _uminus_data_207 = -_cond_data_205;
  wire signed [8-1:0] _cond_data_210;
  assign _cond_data_210 = (__delay_data_761__delay_760_greatereq_208)? _cond_data_205 : _uminus_data_207;
  wire signed [16-1:0] __muladd_madd_odata_211;
  reg signed [16-1:0] __muladd_madd_odata_reg_211;
  wire signed [16-1:0] __muladd_data_211;
  assign __muladd_data_211 = __muladd_madd_odata_reg_211;
  wire __muladd_madd_update_211;
  assign __muladd_madd_update_211 = _mul_9_stream_oready;

  madd_4
  __muladd_madd_211
  (
    .CLK(CLK),
    .update(__muladd_madd_update_211),
    .a(__delay_data_764__delay_763__delay_762__variable_192),
    .b(__delay_data_767__delay_766__delay_765__variable_193),
    .c(_cond_data_210),
    .d(__muladd_madd_odata_211)
  );

  reg [4-1:0] __delay_data_771__delay_770__delay_769____variable_194;
  reg [4-1:0] __delay_data_772__delay_771__delay_770____variable_194;
  reg [4-1:0] __delay_data_773__delay_772__delay_771____variable_194;
  reg [4-1:0] __delay_data_774__delay_773__delay_772____variable_194;
  reg signed [16-1:0] _sra_data_212;
  wire signed [16-1:0] mul_9_z_data;
  assign mul_9_z_data = _sra_data_212;
  wire signed [8-1:0] mul_10_x_data;
  wire signed [8-1:0] mul_10_y_data;
  wire [4-1:0] mul_10_rshift_data;
  reg __mul_10_stream_ivalid_1;
  reg __mul_10_stream_ivalid_2;
  reg __mul_10_stream_ivalid_3;
  reg __mul_10_stream_ivalid_4;
  reg __mul_10_stream_ivalid_5;
  reg __mul_10_stream_ivalid_6;
  reg __mul_10_stream_ivalid_7;
  reg __mul_10_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_216;
  reg [4-1:0] _minus_data_218;
  reg [1-1:0] _greatereq_data_229;
  reg signed [8-1:0] __delay_data_781__variable_213;
  reg signed [8-1:0] __delay_data_784__variable_214;
  reg [4-1:0] __delay_data_787__variable_215;
  reg signed [18-1:0] _sll_data_220;
  reg [1-1:0] __delay_data_778_greaterthan_216;
  reg [1-1:0] __delay_data_779_greatereq_229;
  reg signed [8-1:0] __delay_data_782__delay_781__variable_213;
  reg signed [8-1:0] __delay_data_785__delay_784__variable_214;
  reg [4-1:0] __delay_data_788__delay_787__variable_215;
  reg signed [16-1:0] _cond_data_226;
  reg [1-1:0] __delay_data_780__delay_779_greatereq_229;
  reg signed [8-1:0] __delay_data_783__delay_782__delay_781__variable_213;
  reg signed [8-1:0] __delay_data_786__delay_785__delay_784__variable_214;
  reg [4-1:0] __delay_data_789__delay_788__delay_787__variable_215;
  wire signed [8-1:0] _uminus_data_228;
  assign _uminus_data_228 = -_cond_data_226;
  wire signed [8-1:0] _cond_data_231;
  assign _cond_data_231 = (__delay_data_780__delay_779_greatereq_229)? _cond_data_226 : _uminus_data_228;
  wire signed [16-1:0] __muladd_madd_odata_232;
  reg signed [16-1:0] __muladd_madd_odata_reg_232;
  wire signed [16-1:0] __muladd_data_232;
  assign __muladd_data_232 = __muladd_madd_odata_reg_232;
  wire __muladd_madd_update_232;
  assign __muladd_madd_update_232 = _mul_10_stream_oready;

  madd_5
  __muladd_madd_232
  (
    .CLK(CLK),
    .update(__muladd_madd_update_232),
    .a(__delay_data_783__delay_782__delay_781__variable_213),
    .b(__delay_data_786__delay_785__delay_784__variable_214),
    .c(_cond_data_231),
    .d(__muladd_madd_odata_232)
  );

  reg [4-1:0] __delay_data_790__delay_789__delay_788____variable_215;
  reg [4-1:0] __delay_data_791__delay_790__delay_789____variable_215;
  reg [4-1:0] __delay_data_792__delay_791__delay_790____variable_215;
  reg [4-1:0] __delay_data_793__delay_792__delay_791____variable_215;
  reg signed [16-1:0] _sra_data_233;
  wire signed [16-1:0] mul_10_z_data;
  assign mul_10_z_data = _sra_data_233;
  wire signed [8-1:0] mul_11_x_data;
  wire signed [8-1:0] mul_11_y_data;
  wire [4-1:0] mul_11_rshift_data;
  reg __mul_11_stream_ivalid_1;
  reg __mul_11_stream_ivalid_2;
  reg __mul_11_stream_ivalid_3;
  reg __mul_11_stream_ivalid_4;
  reg __mul_11_stream_ivalid_5;
  reg __mul_11_stream_ivalid_6;
  reg __mul_11_stream_ivalid_7;
  reg __mul_11_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_237;
  reg [4-1:0] _minus_data_239;
  reg [1-1:0] _greatereq_data_250;
  reg signed [8-1:0] __delay_data_800__variable_234;
  reg signed [8-1:0] __delay_data_803__variable_235;
  reg [4-1:0] __delay_data_806__variable_236;
  reg signed [18-1:0] _sll_data_241;
  reg [1-1:0] __delay_data_797_greaterthan_237;
  reg [1-1:0] __delay_data_798_greatereq_250;
  reg signed [8-1:0] __delay_data_801__delay_800__variable_234;
  reg signed [8-1:0] __delay_data_804__delay_803__variable_235;
  reg [4-1:0] __delay_data_807__delay_806__variable_236;
  reg signed [16-1:0] _cond_data_247;
  reg [1-1:0] __delay_data_799__delay_798_greatereq_250;
  reg signed [8-1:0] __delay_data_802__delay_801__delay_800__variable_234;
  reg signed [8-1:0] __delay_data_805__delay_804__delay_803__variable_235;
  reg [4-1:0] __delay_data_808__delay_807__delay_806__variable_236;
  wire signed [8-1:0] _uminus_data_249;
  assign _uminus_data_249 = -_cond_data_247;
  wire signed [8-1:0] _cond_data_252;
  assign _cond_data_252 = (__delay_data_799__delay_798_greatereq_250)? _cond_data_247 : _uminus_data_249;
  wire signed [16-1:0] __muladd_madd_odata_253;
  reg signed [16-1:0] __muladd_madd_odata_reg_253;
  wire signed [16-1:0] __muladd_data_253;
  assign __muladd_data_253 = __muladd_madd_odata_reg_253;
  wire __muladd_madd_update_253;
  assign __muladd_madd_update_253 = _mul_11_stream_oready;

  madd_6
  __muladd_madd_253
  (
    .CLK(CLK),
    .update(__muladd_madd_update_253),
    .a(__delay_data_802__delay_801__delay_800__variable_234),
    .b(__delay_data_805__delay_804__delay_803__variable_235),
    .c(_cond_data_252),
    .d(__muladd_madd_odata_253)
  );

  reg [4-1:0] __delay_data_809__delay_808__delay_807____variable_236;
  reg [4-1:0] __delay_data_810__delay_809__delay_808____variable_236;
  reg [4-1:0] __delay_data_811__delay_810__delay_809____variable_236;
  reg [4-1:0] __delay_data_812__delay_811__delay_810____variable_236;
  reg signed [16-1:0] _sra_data_254;
  wire signed [16-1:0] mul_11_z_data;
  assign mul_11_z_data = _sra_data_254;
  wire signed [8-1:0] mul_12_x_data;
  wire signed [8-1:0] mul_12_y_data;
  wire [4-1:0] mul_12_rshift_data;
  reg __mul_12_stream_ivalid_1;
  reg __mul_12_stream_ivalid_2;
  reg __mul_12_stream_ivalid_3;
  reg __mul_12_stream_ivalid_4;
  reg __mul_12_stream_ivalid_5;
  reg __mul_12_stream_ivalid_6;
  reg __mul_12_stream_ivalid_7;
  reg __mul_12_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_258;
  reg [4-1:0] _minus_data_260;
  reg [1-1:0] _greatereq_data_271;
  reg signed [8-1:0] __delay_data_819__variable_255;
  reg signed [8-1:0] __delay_data_822__variable_256;
  reg [4-1:0] __delay_data_825__variable_257;
  reg signed [18-1:0] _sll_data_262;
  reg [1-1:0] __delay_data_816_greaterthan_258;
  reg [1-1:0] __delay_data_817_greatereq_271;
  reg signed [8-1:0] __delay_data_820__delay_819__variable_255;
  reg signed [8-1:0] __delay_data_823__delay_822__variable_256;
  reg [4-1:0] __delay_data_826__delay_825__variable_257;
  reg signed [16-1:0] _cond_data_268;
  reg [1-1:0] __delay_data_818__delay_817_greatereq_271;
  reg signed [8-1:0] __delay_data_821__delay_820__delay_819__variable_255;
  reg signed [8-1:0] __delay_data_824__delay_823__delay_822__variable_256;
  reg [4-1:0] __delay_data_827__delay_826__delay_825__variable_257;
  wire signed [8-1:0] _uminus_data_270;
  assign _uminus_data_270 = -_cond_data_268;
  wire signed [8-1:0] _cond_data_273;
  assign _cond_data_273 = (__delay_data_818__delay_817_greatereq_271)? _cond_data_268 : _uminus_data_270;
  wire signed [16-1:0] __muladd_madd_odata_274;
  reg signed [16-1:0] __muladd_madd_odata_reg_274;
  wire signed [16-1:0] __muladd_data_274;
  assign __muladd_data_274 = __muladd_madd_odata_reg_274;
  wire __muladd_madd_update_274;
  assign __muladd_madd_update_274 = _mul_12_stream_oready;

  madd_7
  __muladd_madd_274
  (
    .CLK(CLK),
    .update(__muladd_madd_update_274),
    .a(__delay_data_821__delay_820__delay_819__variable_255),
    .b(__delay_data_824__delay_823__delay_822__variable_256),
    .c(_cond_data_273),
    .d(__muladd_madd_odata_274)
  );

  reg [4-1:0] __delay_data_828__delay_827__delay_826____variable_257;
  reg [4-1:0] __delay_data_829__delay_828__delay_827____variable_257;
  reg [4-1:0] __delay_data_830__delay_829__delay_828____variable_257;
  reg [4-1:0] __delay_data_831__delay_830__delay_829____variable_257;
  reg signed [16-1:0] _sra_data_275;
  wire signed [16-1:0] mul_12_z_data;
  assign mul_12_z_data = _sra_data_275;
  wire signed [8-1:0] mul_13_x_data;
  wire signed [8-1:0] mul_13_y_data;
  wire [4-1:0] mul_13_rshift_data;
  reg __mul_13_stream_ivalid_1;
  reg __mul_13_stream_ivalid_2;
  reg __mul_13_stream_ivalid_3;
  reg __mul_13_stream_ivalid_4;
  reg __mul_13_stream_ivalid_5;
  reg __mul_13_stream_ivalid_6;
  reg __mul_13_stream_ivalid_7;
  reg __mul_13_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_279;
  reg [4-1:0] _minus_data_281;
  reg [1-1:0] _greatereq_data_292;
  reg signed [8-1:0] __delay_data_838__variable_276;
  reg signed [8-1:0] __delay_data_841__variable_277;
  reg [4-1:0] __delay_data_844__variable_278;
  reg signed [18-1:0] _sll_data_283;
  reg [1-1:0] __delay_data_835_greaterthan_279;
  reg [1-1:0] __delay_data_836_greatereq_292;
  reg signed [8-1:0] __delay_data_839__delay_838__variable_276;
  reg signed [8-1:0] __delay_data_842__delay_841__variable_277;
  reg [4-1:0] __delay_data_845__delay_844__variable_278;
  reg signed [16-1:0] _cond_data_289;
  reg [1-1:0] __delay_data_837__delay_836_greatereq_292;
  reg signed [8-1:0] __delay_data_840__delay_839__delay_838__variable_276;
  reg signed [8-1:0] __delay_data_843__delay_842__delay_841__variable_277;
  reg [4-1:0] __delay_data_846__delay_845__delay_844__variable_278;
  wire signed [8-1:0] _uminus_data_291;
  assign _uminus_data_291 = -_cond_data_289;
  wire signed [8-1:0] _cond_data_294;
  assign _cond_data_294 = (__delay_data_837__delay_836_greatereq_292)? _cond_data_289 : _uminus_data_291;
  wire signed [16-1:0] __muladd_madd_odata_295;
  reg signed [16-1:0] __muladd_madd_odata_reg_295;
  wire signed [16-1:0] __muladd_data_295;
  assign __muladd_data_295 = __muladd_madd_odata_reg_295;
  wire __muladd_madd_update_295;
  assign __muladd_madd_update_295 = _mul_13_stream_oready;

  madd_8
  __muladd_madd_295
  (
    .CLK(CLK),
    .update(__muladd_madd_update_295),
    .a(__delay_data_840__delay_839__delay_838__variable_276),
    .b(__delay_data_843__delay_842__delay_841__variable_277),
    .c(_cond_data_294),
    .d(__muladd_madd_odata_295)
  );

  reg [4-1:0] __delay_data_847__delay_846__delay_845____variable_278;
  reg [4-1:0] __delay_data_848__delay_847__delay_846____variable_278;
  reg [4-1:0] __delay_data_849__delay_848__delay_847____variable_278;
  reg [4-1:0] __delay_data_850__delay_849__delay_848____variable_278;
  reg signed [16-1:0] _sra_data_296;
  wire signed [16-1:0] mul_13_z_data;
  assign mul_13_z_data = _sra_data_296;
  wire signed [32-1:0] add_tree_3_var0_data;
  wire signed [32-1:0] add_tree_3_var1_data;
  wire signed [32-1:0] add_tree_3_var2_data;
  wire signed [32-1:0] add_tree_3_var3_data;
  wire signed [32-1:0] add_tree_3_var4_data;
  wire signed [32-1:0] add_tree_3_var5_data;
  wire signed [32-1:0] add_tree_3_var6_data;
  wire signed [32-1:0] add_tree_3_var7_data;
  wire signed [32-1:0] add_tree_3_var8_data;
  reg __add_tree_3_stream_ivalid_1;
  reg __add_tree_3_stream_ivalid_2;
  reg signed [32-1:0] __plusn_data_70;
  reg signed [32-1:0] __plusn_data_71;
  reg signed [32-1:0] __plusn_data_72;
  reg signed [32-1:0] __plusn_data_73;
  wire signed [32-1:0] add_tree_3_sum_data;
  assign add_tree_3_sum_data = __plusn_data_73;
  wire signed [32-1:0] acc_1_x_data;
  wire [6-1:0] acc_1_rshift_data;
  wire [32-1:0] acc_1_size_data;
  wire [1-1:0] acc_1__reduce_reset_data;
  reg __acc_1_stream_ivalid_1;
  reg __acc_1_stream_ivalid_2;
  reg __acc_1_stream_ivalid_3;
  reg __acc_1_stream_ivalid_4;
  reg __acc_1_stream_ivalid_5;
  reg [1-1:0] _greaterthan_data_39;
  reg [6-1:0] _minus_data_41;
  reg signed [32-1:0] _reduceadd_data_52;
  reg [33-1:0] _reduceadd_count_52;
  reg _reduceadd_prev_count_max_52;
  wire _reduceadd_reset_cond_52;
  assign _reduceadd_reset_cond_52 = acc_1__reduce_reset_data || _reduceadd_prev_count_max_52;
  wire [33-1:0] _reduceadd_current_count_52;
  assign _reduceadd_current_count_52 = (_reduceadd_reset_cond_52)? 0 : _reduceadd_count_52;
  wire signed [32-1:0] _reduceadd_current_data_52;
  assign _reduceadd_current_data_52 = (_reduceadd_reset_cond_52)? 1'sd0 : _reduceadd_data_52;
  reg [1-1:0] _pulse_data_54;
  reg [33-1:0] _pulse_count_54;
  reg _pulse_prev_count_max_54;
  wire _pulse_reset_cond_54;
  assign _pulse_reset_cond_54 = acc_1__reduce_reset_data || _pulse_prev_count_max_54;
  wire [33-1:0] _pulse_current_count_54;
  assign _pulse_current_count_54 = (_pulse_reset_cond_54)? 0 : _pulse_count_54;
  wire [1-1:0] _pulse_current_data_54;
  assign _pulse_current_data_54 = (_pulse_reset_cond_54)? 1'sd0 : _pulse_data_54;
  reg [6-1:0] __delay_data_859__variable_37;
  reg signed [66-1:0] _sll_data_43;
  reg [1-1:0] __delay_data_856_greaterthan_39;
  reg signed [32-1:0] __delay_data_857_reduceadd_52;
  reg [6-1:0] __delay_data_860__delay_859__variable_37;
  reg [1-1:0] __delay_data_863_pulse_54;
  reg signed [32-1:0] _cond_data_49;
  reg signed [32-1:0] __delay_data_858__delay_857_reduceadd_52;
  reg [6-1:0] __delay_data_861__delay_860__delay_859__variable_37;
  reg [1-1:0] __delay_data_864__delay_863_pulse_54;
  reg signed [32-1:0] _plus_data_56;
  reg [6-1:0] __delay_data_862__delay_861__delay_860__delay_859__variable_37;
  reg [1-1:0] __delay_data_865__delay_864__delay_863_pulse_54;
  reg signed [32-1:0] _sra_data_57;
  reg [1-1:0] __delay_data_866__delay_865__delay_864__delay_863_pulse_54;
  wire signed [32-1:0] acc_1_sum_data;
  assign acc_1_sum_data = _sra_data_57;
  wire [1-1:0] acc_1_valid_data;
  assign acc_1_valid_data = __delay_data_866__delay_865__delay_864__delay_863_pulse_54;
  wire signed [32-1:0] mul_rshift_round_clip_4_x_data;
  wire signed [8-1:0] mul_rshift_round_clip_4_y_data;
  wire [6-1:0] mul_rshift_round_clip_4_rshift_data;
  reg __mul_rshift_round_clip_4_stream_ivalid_1;
  reg __mul_rshift_round_clip_4_stream_ivalid_2;
  reg __mul_rshift_round_clip_4_stream_ivalid_3;
  reg __mul_rshift_round_clip_4_stream_ivalid_4;
  reg __mul_rshift_round_clip_4_stream_ivalid_5;
  reg __mul_rshift_round_clip_4_stream_ivalid_6;
  reg __mul_rshift_round_clip_4_stream_ivalid_7;
  reg __mul_rshift_round_clip_4_stream_ivalid_8;
  wire signed [40-1:0] _times_mul_odata_77;
  reg signed [40-1:0] _times_mul_odata_reg_77;
  wire signed [40-1:0] _times_data_77;
  assign _times_data_77 = _times_mul_odata_reg_77;
  wire _times_mul_update_77;
  assign _times_mul_update_77 = _mul_rshift_round_clip_4_stream_oready;

  multiplier_0
  _times_mul_77
  (
    .CLK(CLK),
    .update(_times_mul_update_77),
    .a(mul_rshift_round_clip_4_x_data),
    .b(mul_rshift_round_clip_4_y_data),
    .c(_times_mul_odata_77)
  );

  wire [6-1:0] _minus_data_80;
  assign _minus_data_80 = mul_rshift_round_clip_4_rshift_data - 2'sd1;
  wire signed [66-1:0] _sll_data_83;
  assign _sll_data_83 = 2'sd1 << _minus_data_80;
  wire [1-1:0] _eq_data_95;
  assign _eq_data_95 = mul_rshift_round_clip_4_rshift_data == 1'sd0;
  reg signed [66-1:0] __delay_data_872_sll_83;
  reg [6-1:0] __delay_data_876__variable_76;
  reg [1-1:0] __delay_data_880_eq_95;
  reg signed [66-1:0] __delay_data_873__delay_872_sll_83;
  reg [6-1:0] __delay_data_877__delay_876__variable_76;
  reg [1-1:0] __delay_data_881__delay_880_eq_95;
  reg signed [66-1:0] __delay_data_874__delay_873__delay_872_sll_83;
  reg [6-1:0] __delay_data_878__delay_877__delay_876__variable_76;
  reg [1-1:0] __delay_data_882__delay_881__delay_880_eq_95;
  reg signed [66-1:0] __delay_data_875__delay_874__delay_873__delay_872_sll_83;
  reg [6-1:0] __delay_data_879__delay_878__delay_877__delay_876__variable_76;
  reg [1-1:0] __delay_data_883__delay_882__delay_881__delay_880_eq_95;
  wire [1-1:0] _pointer_data_78;
  assign _pointer_data_78 = _times_data_77[7'sd39];
  wire signed [2-1:0] _cond_data_90;
  assign _cond_data_90 = (_pointer_data_78)? -2'sd1 : 1'sd0;
  wire signed [41-1:0] _plus_data_91;
  assign _plus_data_91 = _times_data_77 + __delay_data_875__delay_874__delay_873__delay_872_sll_83;
  wire signed [41-1:0] _plus_data_92;
  assign _plus_data_92 = _plus_data_91 + _cond_data_90;
  wire signed [40-1:0] _sra_data_93;
  assign _sra_data_93 = _plus_data_92 >>> __delay_data_879__delay_878__delay_877__delay_876__variable_76;
  reg signed [40-1:0] _cond_data_96;
  reg [1-1:0] _greaterthan_data_97;
  reg [1-1:0] _lessthan_data_101;
  reg [1-1:0] _greatereq_data_105;
  reg signed [40-1:0] __delay_data_884_cond_96;
  reg signed [40-1:0] _cond_data_99;
  reg signed [40-1:0] _cond_data_103;
  reg [1-1:0] __delay_data_885_greatereq_105;
  reg signed [8-1:0] _cond_data_107;
  wire signed [8-1:0] mul_rshift_round_clip_4_z_data;
  assign mul_rshift_round_clip_4_z_data = _cond_data_107;
  reg [33-1:0] _stream_conv2d_24_sink_50_sink_count;
  reg [5-1:0] _stream_conv2d_24_sink_50_sink_mode;
  reg [16-1:0] _stream_conv2d_24_sink_50_sink_generator_id;
  reg [32-1:0] _stream_conv2d_24_sink_50_sink_offset;
  reg [33-1:0] _stream_conv2d_24_sink_50_sink_size;
  reg [32-1:0] _stream_conv2d_24_sink_50_sink_stride;
  reg [32-1:0] _stream_conv2d_24_sink_50_sink_offset_buf;
  reg [33-1:0] _stream_conv2d_24_sink_50_sink_size_buf;
  reg [32-1:0] _stream_conv2d_24_sink_50_sink_stride_buf;
  reg [8-1:0] _stream_conv2d_24_sink_50_sink_sel;
  reg [32-1:0] _stream_conv2d_24_sink_50_sink_waddr;
  reg _stream_conv2d_24_sink_50_sink_wenable;
  reg [8-1:0] _stream_conv2d_24_sink_50_sink_wdata;
  reg _stream_conv2d_24_sink_50_sink_fifo_enq;
  reg [8-1:0] _stream_conv2d_24_sink_50_sink_fifo_wdata;
  reg [8-1:0] _stream_conv2d_24_sink_50_sink_immediate;
  reg [33-1:0] _stream_conv2d_24_sink_51_sink_count;
  reg [5-1:0] _stream_conv2d_24_sink_51_sink_mode;
  reg [16-1:0] _stream_conv2d_24_sink_51_sink_generator_id;
  reg [32-1:0] _stream_conv2d_24_sink_51_sink_offset;
  reg [33-1:0] _stream_conv2d_24_sink_51_sink_size;
  reg [32-1:0] _stream_conv2d_24_sink_51_sink_stride;
  reg [32-1:0] _stream_conv2d_24_sink_51_sink_offset_buf;
  reg [33-1:0] _stream_conv2d_24_sink_51_sink_size_buf;
  reg [32-1:0] _stream_conv2d_24_sink_51_sink_stride_buf;
  reg [8-1:0] _stream_conv2d_24_sink_51_sink_sel;
  reg [32-1:0] _stream_conv2d_24_sink_51_sink_waddr;
  reg _stream_conv2d_24_sink_51_sink_wenable;
  reg [1-1:0] _stream_conv2d_24_sink_51_sink_wdata;
  reg _stream_conv2d_24_sink_51_sink_fifo_enq;
  reg [1-1:0] _stream_conv2d_24_sink_51_sink_fifo_wdata;
  reg [1-1:0] _stream_conv2d_24_sink_51_sink_immediate;
  reg _stream_max_pool_serial_26_stream_ivalid;
  wire _stream_max_pool_serial_26_stream_oready;
  wire _stream_max_pool_serial_26_stream_internal_oready;
  assign _stream_max_pool_serial_26_stream_oready = _stream_max_pool_serial_26_stream_internal_oready;
  reg [32-1:0] _stream_max_pool_serial_26_fsm;
  localparam _stream_max_pool_serial_26_fsm_init = 0;
  wire _stream_max_pool_serial_26_run_flag;
  reg _stream_max_pool_serial_26_source_start;
  wire _stream_max_pool_serial_26_source_stop;
  reg _stream_max_pool_serial_26_source_busy;
  wire _stream_max_pool_serial_26_sink_start;
  wire _stream_max_pool_serial_26_sink_stop;
  wire _stream_max_pool_serial_26_sink_busy;
  wire _stream_max_pool_serial_26_busy;
  reg _stream_max_pool_serial_26_busy_reg;
  wire _stream_max_pool_serial_26_is_root;
  assign _stream_max_pool_serial_26_is_root = 1;
  reg [3-1:0] _stream_max_pool_serial_26_parameter_0_next_parameter_data;
  reg _stream_max_pool_serial_26_source_1_idle;
  reg [33-1:0] _stream_max_pool_serial_26_source_1_source_count;
  reg [5-1:0] _stream_max_pool_serial_26_source_1_source_mode;
  reg [16-1:0] _stream_max_pool_serial_26_source_1_source_generator_id;
  reg [32-1:0] _stream_max_pool_serial_26_source_1_source_offset;
  reg [33-1:0] _stream_max_pool_serial_26_source_1_source_size;
  reg [32-1:0] _stream_max_pool_serial_26_source_1_source_stride;
  reg [32-1:0] _stream_max_pool_serial_26_source_1_source_offset_buf;
  reg [33-1:0] _stream_max_pool_serial_26_source_1_source_size_buf;
  reg [32-1:0] _stream_max_pool_serial_26_source_1_source_stride_buf;
  reg [8-1:0] _stream_max_pool_serial_26_source_1_source_sel;
  reg [32-1:0] _stream_max_pool_serial_26_source_1_source_ram_raddr;
  reg _stream_max_pool_serial_26_source_1_source_ram_renable;
  wire [8-1:0] _stream_max_pool_serial_26_source_1_source_ram_rdata;
  reg _stream_max_pool_serial_26_source_1_source_fifo_deq;
  wire [8-1:0] _stream_max_pool_serial_26_source_1_source_fifo_rdata;
  reg [8-1:0] _stream_max_pool_serial_26_source_1_source_empty_data;
  reg [4-1:0] _stream_max_pool_serial_26_parameter_2_next_parameter_data;
  wire signed [8-1:0] _reduce_max_14_x_data;
  wire [32-1:0] _reduce_max_14_size_data;
  wire [1-1:0] _reduce_max_14__reduce_reset_data;
  reg ___reduce_max_14_stream_ivalid_1;
  reg signed [8-1:0] _reducemax_data_300;
  reg [33-1:0] _reducemax_count_300;
  reg _reducemax_prev_count_max_300;
  wire _reducemax_reset_cond_300;
  assign _reducemax_reset_cond_300 = _reduce_max_14__reduce_reset_data || _reducemax_prev_count_max_300;
  wire [33-1:0] _reducemax_current_count_300;
  assign _reducemax_current_count_300 = (_reducemax_reset_cond_300)? 0 : _reducemax_count_300;
  wire signed [8-1:0] _reducemax_current_data_300;
  assign _reducemax_current_data_300 = (_reducemax_reset_cond_300)? -9'sd128 : _reducemax_data_300;
  reg [1-1:0] _pulse_data_302;
  reg [33-1:0] _pulse_count_302;
  reg _pulse_prev_count_max_302;
  wire _pulse_reset_cond_302;
  assign _pulse_reset_cond_302 = _reduce_max_14__reduce_reset_data || _pulse_prev_count_max_302;
  wire [33-1:0] _pulse_current_count_302;
  assign _pulse_current_count_302 = (_pulse_reset_cond_302)? 0 : _pulse_count_302;
  wire [1-1:0] _pulse_current_data_302;
  assign _pulse_current_data_302 = (_pulse_reset_cond_302)? 1'sd0 : _pulse_data_302;
  wire signed [8-1:0] _reduce_max_14_data_data;
  assign _reduce_max_14_data_data = _reducemax_data_300;
  wire [1-1:0] _reduce_max_14_valid_data;
  assign _reduce_max_14_valid_data = _pulse_data_302;
  reg [33-1:0] _stream_max_pool_serial_26_sink_5_sink_count;
  reg [5-1:0] _stream_max_pool_serial_26_sink_5_sink_mode;
  reg [16-1:0] _stream_max_pool_serial_26_sink_5_sink_generator_id;
  reg [32-1:0] _stream_max_pool_serial_26_sink_5_sink_offset;
  reg [33-1:0] _stream_max_pool_serial_26_sink_5_sink_size;
  reg [32-1:0] _stream_max_pool_serial_26_sink_5_sink_stride;
  reg [32-1:0] _stream_max_pool_serial_26_sink_5_sink_offset_buf;
  reg [33-1:0] _stream_max_pool_serial_26_sink_5_sink_size_buf;
  reg [32-1:0] _stream_max_pool_serial_26_sink_5_sink_stride_buf;
  reg [8-1:0] _stream_max_pool_serial_26_sink_5_sink_sel;
  reg [32-1:0] _stream_max_pool_serial_26_sink_5_sink_waddr;
  reg _stream_max_pool_serial_26_sink_5_sink_wenable;
  reg [8-1:0] _stream_max_pool_serial_26_sink_5_sink_wdata;
  reg _stream_max_pool_serial_26_sink_5_sink_fifo_enq;
  reg [8-1:0] _stream_max_pool_serial_26_sink_5_sink_fifo_wdata;
  reg [8-1:0] _stream_max_pool_serial_26_sink_5_sink_immediate;
  reg [33-1:0] _stream_max_pool_serial_26_sink_6_sink_count;
  reg [5-1:0] _stream_max_pool_serial_26_sink_6_sink_mode;
  reg [16-1:0] _stream_max_pool_serial_26_sink_6_sink_generator_id;
  reg [32-1:0] _stream_max_pool_serial_26_sink_6_sink_offset;
  reg [33-1:0] _stream_max_pool_serial_26_sink_6_sink_size;
  reg [32-1:0] _stream_max_pool_serial_26_sink_6_sink_stride;
  reg [32-1:0] _stream_max_pool_serial_26_sink_6_sink_offset_buf;
  reg [33-1:0] _stream_max_pool_serial_26_sink_6_sink_size_buf;
  reg [32-1:0] _stream_max_pool_serial_26_sink_6_sink_stride_buf;
  reg [8-1:0] _stream_max_pool_serial_26_sink_6_sink_sel;
  reg [32-1:0] _stream_max_pool_serial_26_sink_6_sink_waddr;
  reg _stream_max_pool_serial_26_sink_6_sink_wenable;
  reg [1-1:0] _stream_max_pool_serial_26_sink_6_sink_wdata;
  reg _stream_max_pool_serial_26_sink_6_sink_fifo_enq;
  reg [1-1:0] _stream_max_pool_serial_26_sink_6_sink_fifo_wdata;
  reg [1-1:0] _stream_max_pool_serial_26_sink_6_sink_immediate;
  reg _stream_avg_pool_serial_52_stream_ivalid;
  wire _stream_avg_pool_serial_52_stream_oready;
  wire _stream_avg_pool_serial_52_stream_internal_oready;
  assign _stream_avg_pool_serial_52_stream_oready = _stream_avg_pool_serial_52_stream_internal_oready;
  reg [32-1:0] _stream_avg_pool_serial_52_fsm;
  localparam _stream_avg_pool_serial_52_fsm_init = 0;
  wire _stream_avg_pool_serial_52_run_flag;
  reg _stream_avg_pool_serial_52_source_start;
  wire _stream_avg_pool_serial_52_source_stop;
  reg _stream_avg_pool_serial_52_source_busy;
  wire _stream_avg_pool_serial_52_sink_start;
  wire _stream_avg_pool_serial_52_sink_stop;
  wire _stream_avg_pool_serial_52_sink_busy;
  wire _stream_avg_pool_serial_52_busy;
  reg _stream_avg_pool_serial_52_busy_reg;
  wire _stream_avg_pool_serial_52_is_root;
  assign _stream_avg_pool_serial_52_is_root = 1;
  reg [1-1:0] _stream_avg_pool_serial_52_parameter_0_next_parameter_data;
  reg _stream_avg_pool_serial_52_source_1_idle;
  reg [33-1:0] _stream_avg_pool_serial_52_source_1_source_count;
  reg [5-1:0] _stream_avg_pool_serial_52_source_1_source_mode;
  reg [16-1:0] _stream_avg_pool_serial_52_source_1_source_generator_id;
  reg [32-1:0] _stream_avg_pool_serial_52_source_1_source_offset;
  reg [33-1:0] _stream_avg_pool_serial_52_source_1_source_size;
  reg [32-1:0] _stream_avg_pool_serial_52_source_1_source_stride;
  reg [32-1:0] _stream_avg_pool_serial_52_source_1_source_offset_buf;
  reg [33-1:0] _stream_avg_pool_serial_52_source_1_source_size_buf;
  reg [32-1:0] _stream_avg_pool_serial_52_source_1_source_stride_buf;
  reg [8-1:0] _stream_avg_pool_serial_52_source_1_source_sel;
  reg [32-1:0] _stream_avg_pool_serial_52_source_1_source_ram_raddr;
  reg _stream_avg_pool_serial_52_source_1_source_ram_renable;
  wire [8-1:0] _stream_avg_pool_serial_52_source_1_source_ram_rdata;
  reg _stream_avg_pool_serial_52_source_1_source_fifo_deq;
  wire [8-1:0] _stream_avg_pool_serial_52_source_1_source_fifo_rdata;
  reg [8-1:0] _stream_avg_pool_serial_52_source_1_source_empty_data;
  reg [1-1:0] _stream_avg_pool_serial_52_parameter_2_next_parameter_data;
  wire signed [32-1:0] acc_0_x_data;
  wire [6-1:0] acc_0_rshift_data;
  wire [32-1:0] acc_0_size_data;
  wire [1-1:0] acc_0__reduce_reset_data;
  reg __acc_0_stream_ivalid_1;
  reg __acc_0_stream_ivalid_2;
  reg signed [32-1:0] _reduceadd_data_4;
  reg [33-1:0] _reduceadd_count_4;
  reg _reduceadd_prev_count_max_4;
  wire _reduceadd_reset_cond_4;
  assign _reduceadd_reset_cond_4 = acc_0__reduce_reset_data || _reduceadd_prev_count_max_4;
  wire [33-1:0] _reduceadd_current_count_4;
  assign _reduceadd_current_count_4 = (_reduceadd_reset_cond_4)? 0 : _reduceadd_count_4;
  wire signed [32-1:0] _reduceadd_current_data_4;
  assign _reduceadd_current_data_4 = (_reduceadd_reset_cond_4)? 1'sd0 : _reduceadd_data_4;
  reg [1-1:0] _pulse_data_6;
  reg [33-1:0] _pulse_count_6;
  reg _pulse_prev_count_max_6;
  wire _pulse_reset_cond_6;
  assign _pulse_reset_cond_6 = acc_0__reduce_reset_data || _pulse_prev_count_max_6;
  wire [33-1:0] _pulse_current_count_6;
  assign _pulse_current_count_6 = (_pulse_reset_cond_6)? 0 : _pulse_count_6;
  wire [1-1:0] _pulse_current_data_6;
  assign _pulse_current_data_6 = (_pulse_reset_cond_6)? 1'sd0 : _pulse_data_6;
  wire [5-1:0] _slice_data_12;
  assign _slice_data_12 = acc_0_rshift_data[4'd4:1'd0];
  wire [5-1:0] _minus_data_13;
  assign _minus_data_13 = _slice_data_12 - 2'sd1;
  wire signed [34-1:0] _sll_data_16;
  assign _sll_data_16 = 2'sd1 << _minus_data_13;
  wire [1-1:0] _eq_data_34;
  assign _eq_data_34 = acc_0_rshift_data == 1'sd0;
  reg signed [34-1:0] __delay_data_928_sll_16;
  reg [6-1:0] __delay_data_929__variable_1;
  reg [1-1:0] __delay_data_930_eq_34;
  wire [1-1:0] _pointer_data_8;
  assign _pointer_data_8 = _reduceadd_data_4[6'sd31];
  wire signed [2-1:0] _cond_data_29;
  assign _cond_data_29 = (_pointer_data_8)? -2'sd1 : 1'sd0;
  wire signed [33-1:0] _plus_data_30;
  assign _plus_data_30 = _reduceadd_data_4 + __delay_data_928_sll_16;
  wire signed [33-1:0] _plus_data_31;
  assign _plus_data_31 = _plus_data_30 + _cond_data_29;
  wire signed [32-1:0] _sra_data_32;
  assign _sra_data_32 = _plus_data_31 >>> __delay_data_929__variable_1;
  reg signed [32-1:0] _cond_data_35;
  reg [1-1:0] __delay_data_931_pulse_6;
  wire signed [32-1:0] acc_0_sum_data;
  assign acc_0_sum_data = _cond_data_35;
  wire [1-1:0] acc_0_valid_data;
  assign acc_0_valid_data = __delay_data_931_pulse_6;
  reg [33-1:0] _stream_avg_pool_serial_52_sink_5_sink_count;
  reg [5-1:0] _stream_avg_pool_serial_52_sink_5_sink_mode;
  reg [16-1:0] _stream_avg_pool_serial_52_sink_5_sink_generator_id;
  reg [32-1:0] _stream_avg_pool_serial_52_sink_5_sink_offset;
  reg [33-1:0] _stream_avg_pool_serial_52_sink_5_sink_size;
  reg [32-1:0] _stream_avg_pool_serial_52_sink_5_sink_stride;
  reg [32-1:0] _stream_avg_pool_serial_52_sink_5_sink_offset_buf;
  reg [33-1:0] _stream_avg_pool_serial_52_sink_5_sink_size_buf;
  reg [32-1:0] _stream_avg_pool_serial_52_sink_5_sink_stride_buf;
  reg [8-1:0] _stream_avg_pool_serial_52_sink_5_sink_sel;
  reg [32-1:0] _stream_avg_pool_serial_52_sink_5_sink_waddr;
  reg _stream_avg_pool_serial_52_sink_5_sink_wenable;
  reg [8-1:0] _stream_avg_pool_serial_52_sink_5_sink_wdata;
  reg _stream_avg_pool_serial_52_sink_5_sink_fifo_enq;
  reg [8-1:0] _stream_avg_pool_serial_52_sink_5_sink_fifo_wdata;
  reg [8-1:0] _stream_avg_pool_serial_52_sink_5_sink_immediate;
  reg [33-1:0] _stream_avg_pool_serial_52_sink_6_sink_count;
  reg [5-1:0] _stream_avg_pool_serial_52_sink_6_sink_mode;
  reg [16-1:0] _stream_avg_pool_serial_52_sink_6_sink_generator_id;
  reg [32-1:0] _stream_avg_pool_serial_52_sink_6_sink_offset;
  reg [33-1:0] _stream_avg_pool_serial_52_sink_6_sink_size;
  reg [32-1:0] _stream_avg_pool_serial_52_sink_6_sink_stride;
  reg [32-1:0] _stream_avg_pool_serial_52_sink_6_sink_offset_buf;
  reg [33-1:0] _stream_avg_pool_serial_52_sink_6_sink_size_buf;
  reg [32-1:0] _stream_avg_pool_serial_52_sink_6_sink_stride_buf;
  reg [8-1:0] _stream_avg_pool_serial_52_sink_6_sink_sel;
  reg [32-1:0] _stream_avg_pool_serial_52_sink_6_sink_waddr;
  reg _stream_avg_pool_serial_52_sink_6_sink_wenable;
  reg [1-1:0] _stream_avg_pool_serial_52_sink_6_sink_wdata;
  reg _stream_avg_pool_serial_52_sink_6_sink_fifo_enq;
  reg [1-1:0] _stream_avg_pool_serial_52_sink_6_sink_fifo_wdata;
  reg [1-1:0] _stream_avg_pool_serial_52_sink_6_sink_immediate;
  reg _stream_matmul_55_stream_ivalid;
  wire _stream_matmul_55_stream_oready;
  wire _stream_matmul_55_stream_internal_oready;
  assign _stream_matmul_55_stream_oready = _stream_matmul_55_stream_internal_oready;
  reg [32-1:0] _stream_matmul_55_fsm;
  localparam _stream_matmul_55_fsm_init = 0;
  wire _stream_matmul_55_run_flag;
  reg _stream_matmul_55_source_start;
  wire _stream_matmul_55_source_stop;
  reg _stream_matmul_55_source_busy;
  wire _stream_matmul_55_sink_start;
  wire _stream_matmul_55_sink_stop;
  wire _stream_matmul_55_sink_busy;
  wire _stream_matmul_55_busy;
  reg _stream_matmul_55_busy_reg;
  wire _stream_matmul_55_is_root;
  assign _stream_matmul_55_is_root = 1;
  reg [15-1:0] _stream_matmul_55_parameter_0_next_parameter_data;
  reg [1-1:0] _stream_matmul_55_parameter_1_next_parameter_data;
  reg [1-1:0] _stream_matmul_55_parameter_2_next_parameter_data;
  reg [1-1:0] _stream_matmul_55_parameter_3_next_parameter_data;
  reg [1-1:0] _stream_matmul_55_parameter_4_next_parameter_data;
  reg [1-1:0] _stream_matmul_55_parameter_6_next_parameter_data;
  reg _stream_matmul_55_source_7_idle;
  reg [33-1:0] _stream_matmul_55_source_7_source_count;
  reg [5-1:0] _stream_matmul_55_source_7_source_mode;
  reg [16-1:0] _stream_matmul_55_source_7_source_generator_id;
  reg [32-1:0] _stream_matmul_55_source_7_source_offset;
  reg [33-1:0] _stream_matmul_55_source_7_source_size;
  reg [32-1:0] _stream_matmul_55_source_7_source_stride;
  reg [32-1:0] _stream_matmul_55_source_7_source_offset_buf;
  reg [33-1:0] _stream_matmul_55_source_7_source_size_buf;
  reg [32-1:0] _stream_matmul_55_source_7_source_stride_buf;
  reg [8-1:0] _stream_matmul_55_source_7_source_sel;
  reg [32-1:0] _stream_matmul_55_source_7_source_ram_raddr;
  reg _stream_matmul_55_source_7_source_ram_renable;
  wire [32-1:0] _stream_matmul_55_source_7_source_ram_rdata;
  reg _stream_matmul_55_source_7_source_fifo_deq;
  wire [32-1:0] _stream_matmul_55_source_7_source_fifo_rdata;
  reg [32-1:0] _stream_matmul_55_source_7_source_empty_data;
  reg [1-1:0] _stream_matmul_55_parameter_8_next_parameter_data;
  reg _stream_matmul_55_source_9_idle;
  reg [33-1:0] _stream_matmul_55_source_9_source_count;
  reg [5-1:0] _stream_matmul_55_source_9_source_mode;
  reg [16-1:0] _stream_matmul_55_source_9_source_generator_id;
  reg [32-1:0] _stream_matmul_55_source_9_source_offset;
  reg [33-1:0] _stream_matmul_55_source_9_source_size;
  reg [32-1:0] _stream_matmul_55_source_9_source_stride;
  reg [32-1:0] _stream_matmul_55_source_9_source_offset_buf;
  reg [33-1:0] _stream_matmul_55_source_9_source_size_buf;
  reg [32-1:0] _stream_matmul_55_source_9_source_stride_buf;
  reg [8-1:0] _stream_matmul_55_source_9_source_sel;
  reg [32-1:0] _stream_matmul_55_source_9_source_ram_raddr;
  reg _stream_matmul_55_source_9_source_ram_renable;
  wire [8-1:0] _stream_matmul_55_source_9_source_ram_rdata;
  reg _stream_matmul_55_source_9_source_fifo_deq;
  wire [8-1:0] _stream_matmul_55_source_9_source_fifo_rdata;
  reg [8-1:0] _stream_matmul_55_source_9_source_empty_data;
  reg [1-1:0] _stream_matmul_55_parameter_10_next_parameter_data;
  reg _stream_matmul_55_source_11_idle;
  reg [33-1:0] _stream_matmul_55_source_11_source_count;
  reg [5-1:0] _stream_matmul_55_source_11_source_mode;
  reg [16-1:0] _stream_matmul_55_source_11_source_generator_id;
  reg [32-1:0] _stream_matmul_55_source_11_source_offset;
  reg [33-1:0] _stream_matmul_55_source_11_source_size;
  reg [32-1:0] _stream_matmul_55_source_11_source_stride;
  reg [32-1:0] _stream_matmul_55_source_11_source_offset_buf;
  reg [33-1:0] _stream_matmul_55_source_11_source_size_buf;
  reg [32-1:0] _stream_matmul_55_source_11_source_stride_buf;
  reg [8-1:0] _stream_matmul_55_source_11_source_sel;
  reg [32-1:0] _stream_matmul_55_source_11_source_ram_raddr;
  reg _stream_matmul_55_source_11_source_ram_renable;
  wire [8-1:0] _stream_matmul_55_source_11_source_ram_rdata;
  reg _stream_matmul_55_source_11_source_fifo_deq;
  wire [8-1:0] _stream_matmul_55_source_11_source_fifo_rdata;
  reg [8-1:0] _stream_matmul_55_source_11_source_empty_data;
  reg [1-1:0] _stream_matmul_55_parameter_12_next_parameter_data;
  reg _stream_matmul_55_source_13_idle;
  reg [33-1:0] _stream_matmul_55_source_13_source_count;
  reg [5-1:0] _stream_matmul_55_source_13_source_mode;
  reg [16-1:0] _stream_matmul_55_source_13_source_generator_id;
  reg [32-1:0] _stream_matmul_55_source_13_source_offset;
  reg [33-1:0] _stream_matmul_55_source_13_source_size;
  reg [32-1:0] _stream_matmul_55_source_13_source_stride;
  reg [32-1:0] _stream_matmul_55_source_13_source_offset_buf;
  reg [33-1:0] _stream_matmul_55_source_13_source_size_buf;
  reg [32-1:0] _stream_matmul_55_source_13_source_stride_buf;
  reg [8-1:0] _stream_matmul_55_source_13_source_sel;
  reg [32-1:0] _stream_matmul_55_source_13_source_ram_raddr;
  reg _stream_matmul_55_source_13_source_ram_renable;
  wire [8-1:0] _stream_matmul_55_source_13_source_ram_rdata;
  reg _stream_matmul_55_source_13_source_fifo_deq;
  wire [8-1:0] _stream_matmul_55_source_13_source_fifo_rdata;
  reg [8-1:0] _stream_matmul_55_source_13_source_empty_data;
  reg [1-1:0] _stream_matmul_55_parameter_14_next_parameter_data;
  reg _stream_matmul_55_source_15_idle;
  reg [33-1:0] _stream_matmul_55_source_15_source_count;
  reg [5-1:0] _stream_matmul_55_source_15_source_mode;
  reg [16-1:0] _stream_matmul_55_source_15_source_generator_id;
  reg [32-1:0] _stream_matmul_55_source_15_source_offset;
  reg [33-1:0] _stream_matmul_55_source_15_source_size;
  reg [32-1:0] _stream_matmul_55_source_15_source_stride;
  reg [32-1:0] _stream_matmul_55_source_15_source_offset_buf;
  reg [33-1:0] _stream_matmul_55_source_15_source_size_buf;
  reg [32-1:0] _stream_matmul_55_source_15_source_stride_buf;
  reg [8-1:0] _stream_matmul_55_source_15_source_sel;
  reg [32-1:0] _stream_matmul_55_source_15_source_ram_raddr;
  reg _stream_matmul_55_source_15_source_ram_renable;
  wire [8-1:0] _stream_matmul_55_source_15_source_ram_rdata;
  reg _stream_matmul_55_source_15_source_fifo_deq;
  wire [8-1:0] _stream_matmul_55_source_15_source_fifo_rdata;
  reg [8-1:0] _stream_matmul_55_source_15_source_empty_data;
  reg [1-1:0] _stream_matmul_55_parameter_16_next_parameter_data;
  reg [1-1:0] _stream_matmul_55_parameter_17_next_parameter_data;
  reg [5-1:0] _stream_matmul_55_parameter_18_next_parameter_data;
  reg [2-1:0] _stream_matmul_55_parameter_19_next_parameter_data;
  reg _stream_matmul_55_source_20_idle;
  reg [33-1:0] _stream_matmul_55_source_20_source_count;
  reg [5-1:0] _stream_matmul_55_source_20_source_mode;
  reg [16-1:0] _stream_matmul_55_source_20_source_generator_id;
  reg [32-1:0] _stream_matmul_55_source_20_source_offset;
  reg [33-1:0] _stream_matmul_55_source_20_source_size;
  reg [32-1:0] _stream_matmul_55_source_20_source_stride;
  reg [32-1:0] _stream_matmul_55_source_20_source_offset_buf;
  reg [33-1:0] _stream_matmul_55_source_20_source_size_buf;
  reg [32-1:0] _stream_matmul_55_source_20_source_stride_buf;
  reg [8-1:0] _stream_matmul_55_source_20_source_sel;
  reg [32-1:0] _stream_matmul_55_source_20_source_ram_raddr;
  reg _stream_matmul_55_source_20_source_ram_renable;
  wire [8-1:0] _stream_matmul_55_source_20_source_ram_rdata;
  reg _stream_matmul_55_source_20_source_fifo_deq;
  wire [8-1:0] _stream_matmul_55_source_20_source_fifo_rdata;
  reg [8-1:0] _stream_matmul_55_source_20_source_empty_data;
  reg _stream_matmul_55_source_21_idle;
  reg [33-1:0] _stream_matmul_55_source_21_source_count;
  reg [5-1:0] _stream_matmul_55_source_21_source_mode;
  reg [16-1:0] _stream_matmul_55_source_21_source_generator_id;
  reg [32-1:0] _stream_matmul_55_source_21_source_offset;
  reg [33-1:0] _stream_matmul_55_source_21_source_size;
  reg [32-1:0] _stream_matmul_55_source_21_source_stride;
  reg [32-1:0] _stream_matmul_55_source_21_source_offset_buf;
  reg [33-1:0] _stream_matmul_55_source_21_source_size_buf;
  reg [32-1:0] _stream_matmul_55_source_21_source_stride_buf;
  reg [8-1:0] _stream_matmul_55_source_21_source_sel;
  reg [32-1:0] _stream_matmul_55_source_21_source_ram_raddr;
  reg _stream_matmul_55_source_21_source_ram_renable;
  wire [8-1:0] _stream_matmul_55_source_21_source_ram_rdata;
  reg _stream_matmul_55_source_21_source_fifo_deq;
  wire [8-1:0] _stream_matmul_55_source_21_source_fifo_rdata;
  reg [8-1:0] _stream_matmul_55_source_21_source_empty_data;
  wire signed [32-1:0] add_tree_2_var0_data;
  wire signed [32-1:0] _cast_src_59;
  assign _cast_src_59 = add_tree_2_var0_data;
  wire signed [32-1:0] _cast_data_59;
  assign _cast_data_59 = _cast_src_59;
  wire signed [32-1:0] add_tree_2_sum_data;
  assign add_tree_2_sum_data = _cast_data_59;
  reg [33-1:0] _stream_matmul_55_sink_26_sink_count;
  reg [5-1:0] _stream_matmul_55_sink_26_sink_mode;
  reg [16-1:0] _stream_matmul_55_sink_26_sink_generator_id;
  reg [32-1:0] _stream_matmul_55_sink_26_sink_offset;
  reg [33-1:0] _stream_matmul_55_sink_26_sink_size;
  reg [32-1:0] _stream_matmul_55_sink_26_sink_stride;
  reg [32-1:0] _stream_matmul_55_sink_26_sink_offset_buf;
  reg [33-1:0] _stream_matmul_55_sink_26_sink_size_buf;
  reg [32-1:0] _stream_matmul_55_sink_26_sink_stride_buf;
  reg [8-1:0] _stream_matmul_55_sink_26_sink_sel;
  reg [32-1:0] _stream_matmul_55_sink_26_sink_waddr;
  reg _stream_matmul_55_sink_26_sink_wenable;
  reg [8-1:0] _stream_matmul_55_sink_26_sink_wdata;
  reg _stream_matmul_55_sink_26_sink_fifo_enq;
  reg [8-1:0] _stream_matmul_55_sink_26_sink_fifo_wdata;
  reg [8-1:0] _stream_matmul_55_sink_26_sink_immediate;
  reg [33-1:0] _stream_matmul_55_sink_27_sink_count;
  reg [5-1:0] _stream_matmul_55_sink_27_sink_mode;
  reg [16-1:0] _stream_matmul_55_sink_27_sink_generator_id;
  reg [32-1:0] _stream_matmul_55_sink_27_sink_offset;
  reg [33-1:0] _stream_matmul_55_sink_27_sink_size;
  reg [32-1:0] _stream_matmul_55_sink_27_sink_stride;
  reg [32-1:0] _stream_matmul_55_sink_27_sink_offset_buf;
  reg [33-1:0] _stream_matmul_55_sink_27_sink_size_buf;
  reg [32-1:0] _stream_matmul_55_sink_27_sink_stride_buf;
  reg [8-1:0] _stream_matmul_55_sink_27_sink_sel;
  reg [32-1:0] _stream_matmul_55_sink_27_sink_waddr;
  reg _stream_matmul_55_sink_27_sink_wenable;
  reg [1-1:0] _stream_matmul_55_sink_27_sink_wdata;
  reg _stream_matmul_55_sink_27_sink_fifo_enq;
  reg [1-1:0] _stream_matmul_55_sink_27_sink_fifo_wdata;
  reg [1-1:0] _stream_matmul_55_sink_27_sink_immediate;
  reg [32-1:0] main_fsm;
  localparam main_fsm_init = 0;
  reg [32-1:0] internal_state_counter;
  reg [32-1:0] conv2d_24_objaddr;
  reg [32-1:0] conv2d_24_arg_objaddr_0;
  reg [32-1:0] conv2d_24_arg_objaddr_1;
  reg [32-1:0] conv2d_24_arg_objaddr_2;
  reg [32-1:0] conv2d_24_arg_objaddr_3;
  reg [32-1:0] control_conv2d_24;
  localparam control_conv2d_24_init = 0;
  reg _control_conv2d_24_called;
  wire signed [32-1:0] conv2d_24_act_base_offset;
  reg signed [32-1:0] conv2d_24_act_base_offset_row;
  reg signed [32-1:0] conv2d_24_act_base_offset_bat;
  assign conv2d_24_act_base_offset = conv2d_24_act_base_offset_row + conv2d_24_act_base_offset_bat;
  reg signed [32-1:0] conv2d_24_filter_base_offset;
  reg [32-1:0] conv2d_24_next_stream_num_ops;
  wire signed [32-1:0] conv2d_24_out_base_offset;
  reg signed [32-1:0] conv2d_24_out_base_offset_val;
  reg signed [32-1:0] conv2d_24_out_base_offset_col;
  reg signed [32-1:0] conv2d_24_out_base_offset_row;
  reg signed [32-1:0] conv2d_24_out_base_offset_bat;
  reg signed [32-1:0] conv2d_24_out_base_offset_och;
  assign conv2d_24_out_base_offset = conv2d_24_out_base_offset_val + conv2d_24_out_base_offset_col + conv2d_24_out_base_offset_row + conv2d_24_out_base_offset_bat + conv2d_24_out_base_offset_och;
  reg conv2d_24_dma_flag_0;
  reg conv2d_24_dma_flag_1;
  reg conv2d_24_dma_flag_2;
  reg [32-1:0] conv2d_24_sync_comp_count;
  reg [32-1:0] conv2d_24_sync_out_count;
  reg [32-1:0] conv2d_24_write_count;
  reg [32-1:0] conv2d_24_next_out_write_size;
  reg [32-1:0] conv2d_24_col_count;
  reg [32-1:0] conv2d_24_row_count;
  reg [32-1:0] conv2d_24_bat_count;
  reg [32-1:0] conv2d_24_och_count;
  reg [2-1:0] conv2d_24_col_select;
  reg [2-1:0] conv2d_24_row_select;
  reg [32-1:0] conv2d_24_out_col_count;
  reg [32-1:0] conv2d_24_out_row_count;
  reg [32-1:0] conv2d_24_out_ram_select;
  reg [32-1:0] conv2d_24_prev_col_count;
  reg [32-1:0] conv2d_24_prev_row_count;
  reg [32-1:0] conv2d_24_prev_bat_count;
  reg [32-1:0] conv2d_24_prev_och_count;
  reg [2-1:0] conv2d_24_prev_row_select;
  reg [32-1:0] conv2d_24_stream_act_local_0;
  reg [32-1:0] conv2d_24_stream_act_local_1;
  reg [32-1:0] conv2d_24_stream_act_local_2;
  reg [32-1:0] conv2d_24_stream_act_local_3;
  reg [32-1:0] conv2d_24_stream_act_local_4;
  reg [32-1:0] conv2d_24_stream_act_local_5;
  reg [32-1:0] conv2d_24_stream_act_local_6;
  reg [32-1:0] conv2d_24_stream_act_local_7;
  reg [32-1:0] conv2d_24_stream_act_local_8;
  reg [32-1:0] conv2d_24_stream_out_local_val;
  reg [32-1:0] conv2d_24_stream_out_local_col;
  wire [32-1:0] conv2d_24_stream_out_local;
  assign conv2d_24_stream_out_local = conv2d_24_stream_out_local_val + conv2d_24_stream_out_local_col;
  reg [32-1:0] conv2d_24_act_page_comp_offset_0;
  reg [32-1:0] conv2d_24_act_page_comp_offset_1;
  reg [32-1:0] conv2d_24_act_page_comp_offset_2;
  reg [32-1:0] conv2d_24_act_page_dma_offset_0;
  reg [32-1:0] conv2d_24_act_page_dma_offset_1;
  reg [32-1:0] conv2d_24_act_page_dma_offset_2;
  reg [32-1:0] conv2d_24_filter_page_comp_offset;
  reg [32-1:0] conv2d_24_filter_page_dma_offset;
  reg conv2d_24_out_page;
  reg [32-1:0] conv2d_24_out_page_comp_offset;
  reg [32-1:0] conv2d_24_out_page_dma_offset;
  reg [32-1:0] conv2d_24_out_laddr_offset;
  reg conv2d_24_skip_read_filter;
  reg conv2d_24_skip_read_act;
  reg conv2d_24_skip_comp;
  reg conv2d_24_skip_write_out;
  wire [32-1:0] mask_addr_shifted_54;
  assign mask_addr_shifted_54 = conv2d_24_arg_objaddr_2 + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_55;
  assign mask_addr_masked_55 = mask_addr_shifted_54 << 2;
  reg [32-1:0] _maxi_read_req_fsm;
  localparam _maxi_read_req_fsm_init = 0;
  reg [33-1:0] _maxi_read_cur_global_size;
  reg _maxi_read_cont;
  wire [8-1:0] pack_read_req_op_sel_56;
  wire [32-1:0] pack_read_req_local_addr_57;
  wire [32-1:0] pack_read_req_local_stride_58;
  wire [33-1:0] pack_read_req_local_size_59;
  wire [32-1:0] pack_read_req_local_blocksize_60;
  assign pack_read_req_op_sel_56 = _maxi_read_op_sel;
  assign pack_read_req_local_addr_57 = _maxi_read_local_addr;
  assign pack_read_req_local_stride_58 = _maxi_read_local_stride;
  assign pack_read_req_local_size_59 = _maxi_read_local_size;
  assign pack_read_req_local_blocksize_60 = _maxi_read_local_blocksize;
  wire [137-1:0] pack_read_req_packed_61;
  assign pack_read_req_packed_61 = { pack_read_req_op_sel_56, pack_read_req_local_addr_57, pack_read_req_local_stride_58, pack_read_req_local_size_59, pack_read_req_local_blocksize_60 };
  assign _maxi_read_req_fifo_wdata = ((_maxi_read_req_fsm == 0) && _maxi_read_start && !_maxi_read_req_fifo_almost_full)? pack_read_req_packed_61 : 'hx;
  assign _maxi_read_req_fifo_enq = ((_maxi_read_req_fsm == 0) && _maxi_read_start && !_maxi_read_req_fifo_almost_full)? (_maxi_read_req_fsm == 0) && _maxi_read_start && !_maxi_read_req_fifo_almost_full && !_maxi_read_req_fifo_almost_full : 0;
  localparam _tmp_62 = 1;
  wire [_tmp_62-1:0] _tmp_63;
  assign _tmp_63 = !_maxi_read_req_fifo_almost_full;
  reg [_tmp_62-1:0] __tmp_63_1;
  wire [32-1:0] mask_addr_shifted_64;
  assign mask_addr_shifted_64 = _maxi_read_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_65;
  assign mask_addr_masked_65 = mask_addr_shifted_64 << 2;
  wire [32-1:0] mask_addr_shifted_66;
  assign mask_addr_shifted_66 = _maxi_read_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_67;
  assign mask_addr_masked_67 = mask_addr_shifted_66 << 2;
  wire [32-1:0] mask_addr_shifted_68;
  assign mask_addr_shifted_68 = _maxi_read_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_69;
  assign mask_addr_masked_69 = mask_addr_shifted_68 << 2;
  wire [32-1:0] mask_addr_shifted_70;
  assign mask_addr_shifted_70 = _maxi_read_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_71;
  assign mask_addr_masked_71 = mask_addr_shifted_70 << 2;
  wire [32-1:0] mask_addr_shifted_72;
  assign mask_addr_shifted_72 = _maxi_read_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_73;
  assign mask_addr_masked_73 = mask_addr_shifted_72 << 2;
  wire [32-1:0] mask_addr_shifted_74;
  assign mask_addr_shifted_74 = _maxi_read_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_75;
  assign mask_addr_masked_75 = mask_addr_shifted_74 << 2;
  reg _maxi_raddr_cond_0_1;
  reg [32-1:0] _maxi_read_data_fsm;
  localparam _maxi_read_data_fsm_init = 0;
  reg [32-1:0] write_burst_fsm_0;
  localparam write_burst_fsm_0_init = 0;
  reg [12-1:0] write_burst_addr_76;
  reg [12-1:0] write_burst_stride_77;
  reg [33-1:0] write_burst_length_78;
  reg write_burst_done_79;
  assign ram_w32_l4096_id0_1_addr = ((write_burst_fsm_0 == 1) && _maxi_rvalid_sb_0)? write_burst_addr_76 : 'hx;
  assign ram_w32_l4096_id0_1_wdata = ((write_burst_fsm_0 == 1) && _maxi_rvalid_sb_0)? _maxi_rdata_sb_0 : 'hx;
  assign ram_w32_l4096_id0_1_wenable = ((write_burst_fsm_0 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  assign ram_w32_l4096_id0_1_enable = ((write_burst_fsm_0 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  wire [1-1:0] _dma_read_packed_high_local_size_80;
  assign _dma_read_packed_high_local_size_80 = cparam_conv2d_24_scale_num >> 2;
  wire [2-1:0] _dma_read_packed_low_local_size_81;
  assign _dma_read_packed_low_local_size_81 = cparam_conv2d_24_scale_num & { 2{ 1'd1 } };
  wire [1-1:0] _dma_read_packed_local_packed_size_82;
  assign _dma_read_packed_local_packed_size_82 = (_dma_read_packed_low_local_size_81 > 0)? _dma_read_packed_high_local_size_80 + 1 : _dma_read_packed_high_local_size_80;
  wire [32-1:0] mask_addr_shifted_83;
  assign mask_addr_shifted_83 = conv2d_24_arg_objaddr_3 + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_84;
  assign mask_addr_masked_84 = mask_addr_shifted_83 << 2;
  reg [32-1:0] write_burst_packed_fsm_1;
  localparam write_burst_packed_fsm_1_init = 0;
  reg [11-1:0] write_burst_packed_addr_85;
  reg [11-1:0] write_burst_packed_stride_86;
  reg [33-1:0] write_burst_packed_length_87;
  reg write_burst_packed_done_88;
  wire [9-1:0] write_burst_packed_ram_addr_89;
  assign write_burst_packed_ram_addr_89 = write_burst_packed_addr_85 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_90;
  assign write_burst_packed_ram_wdata_90 = _maxi_rdata_sb_0 >> 0;
  assign ram_w8_l2048_id0_0_1_addr = ((write_burst_packed_fsm_1 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_addr_89 : 'hx;
  assign ram_w8_l2048_id0_0_1_wdata = ((write_burst_packed_fsm_1 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_wdata_90 : 'hx;
  assign ram_w8_l2048_id0_0_1_wenable = ((write_burst_packed_fsm_1 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  assign ram_w8_l2048_id0_0_1_enable = ((write_burst_packed_fsm_1 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  wire [9-1:0] write_burst_packed_ram_addr_91;
  assign write_burst_packed_ram_addr_91 = write_burst_packed_addr_85 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_92;
  assign write_burst_packed_ram_wdata_92 = _maxi_rdata_sb_0 >> 8;
  assign ram_w8_l2048_id0_1_1_addr = ((write_burst_packed_fsm_1 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_addr_91 : 'hx;
  assign ram_w8_l2048_id0_1_1_wdata = ((write_burst_packed_fsm_1 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_wdata_92 : 'hx;
  assign ram_w8_l2048_id0_1_1_wenable = ((write_burst_packed_fsm_1 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  assign ram_w8_l2048_id0_1_1_enable = ((write_burst_packed_fsm_1 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  wire [9-1:0] write_burst_packed_ram_addr_93;
  assign write_burst_packed_ram_addr_93 = write_burst_packed_addr_85 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_94;
  assign write_burst_packed_ram_wdata_94 = _maxi_rdata_sb_0 >> 16;
  assign ram_w8_l2048_id0_2_1_addr = ((write_burst_packed_fsm_1 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_addr_93 : 'hx;
  assign ram_w8_l2048_id0_2_1_wdata = ((write_burst_packed_fsm_1 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_wdata_94 : 'hx;
  assign ram_w8_l2048_id0_2_1_wenable = ((write_burst_packed_fsm_1 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  assign ram_w8_l2048_id0_2_1_enable = ((write_burst_packed_fsm_1 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  wire [9-1:0] write_burst_packed_ram_addr_95;
  assign write_burst_packed_ram_addr_95 = write_burst_packed_addr_85 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_96;
  assign write_burst_packed_ram_wdata_96 = _maxi_rdata_sb_0 >> 24;
  assign ram_w8_l2048_id0_3_1_addr = ((write_burst_packed_fsm_1 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_addr_95 : 'hx;
  assign ram_w8_l2048_id0_3_1_wdata = ((write_burst_packed_fsm_1 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_wdata_96 : 'hx;
  assign ram_w8_l2048_id0_3_1_wenable = ((write_burst_packed_fsm_1 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  assign ram_w8_l2048_id0_3_1_enable = ((write_burst_packed_fsm_1 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  wire [15-1:0] _dma_write_block_high_local_size_97;
  assign _dma_write_block_high_local_size_97 = cparam_conv2d_24_filter_read_size >> 2;
  wire [2-1:0] _dma_write_block_low_local_size_98;
  assign _dma_write_block_low_local_size_98 = cparam_conv2d_24_filter_read_size & { 2{ 1'd1 } };
  wire [15-1:0] _dma_write_block_local_size_99;
  assign _dma_write_block_local_size_99 = (_dma_write_block_low_local_size_98 > 0)? _dma_write_block_high_local_size_97 + 1 : _dma_write_block_high_local_size_97;
  wire [10-1:0] _dma_read_block_high_local_blocksize_100;
  assign _dma_read_block_high_local_blocksize_100 = cparam_conv2d_24_filter_read_block >> 2;
  wire [3-1:0] _dma_read_block_low_local_blocksize_101;
  assign _dma_read_block_low_local_blocksize_101 = cparam_conv2d_24_filter_read_block & { 2{ 1'd1 } };
  wire [10-1:0] _dma_read_block_local_blocksize_102;
  assign _dma_read_block_local_blocksize_102 = (_dma_read_block_low_local_blocksize_101 > 0)? _dma_read_block_high_local_blocksize_100 + 1 : _dma_read_block_high_local_blocksize_100;
  wire [32-1:0] mask_addr_shifted_103;
  assign mask_addr_shifted_103 = conv2d_24_arg_objaddr_1 + conv2d_24_filter_base_offset + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_104;
  assign mask_addr_masked_104 = mask_addr_shifted_103 << 2;
  wire write_burst_block_ram_wvalid_105;
  wire write_burst_block_ram_wquit_106;
  reg [32-1:0] write_burst_packed_fsm_2;
  localparam write_burst_packed_fsm_2_init = 0;
  reg [12-1:0] write_burst_packed_addr_107;
  reg [12-1:0] write_burst_packed_stride_108;
  reg [33-1:0] write_burst_packed_length_109;
  reg write_burst_packed_done_110;
  wire [10-1:0] write_burst_packed_ram_addr_111;
  assign write_burst_packed_ram_addr_111 = write_burst_packed_addr_107 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_112;
  assign write_burst_packed_ram_wdata_112 = _maxi_rdata_sb_0 >> 0;
  assign ram_w8_l4096_id0_0_1_addr = ((write_burst_packed_fsm_2 == 1) && write_burst_block_ram_wvalid_105)? write_burst_packed_ram_addr_111 : 'hx;
  assign ram_w8_l4096_id0_0_1_wdata = ((write_burst_packed_fsm_2 == 1) && write_burst_block_ram_wvalid_105)? write_burst_packed_ram_wdata_112 : 'hx;
  assign ram_w8_l4096_id0_0_1_wenable = ((write_burst_packed_fsm_2 == 1) && write_burst_block_ram_wvalid_105)? 1'd1 : 0;
  assign ram_w8_l4096_id0_0_1_enable = ((write_burst_packed_fsm_2 == 1) && write_burst_block_ram_wvalid_105)? 1'd1 : 0;
  wire [10-1:0] write_burst_packed_ram_addr_113;
  assign write_burst_packed_ram_addr_113 = write_burst_packed_addr_107 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_114;
  assign write_burst_packed_ram_wdata_114 = _maxi_rdata_sb_0 >> 8;
  assign ram_w8_l4096_id0_1_1_addr = ((write_burst_packed_fsm_2 == 1) && write_burst_block_ram_wvalid_105)? write_burst_packed_ram_addr_113 : 'hx;
  assign ram_w8_l4096_id0_1_1_wdata = ((write_burst_packed_fsm_2 == 1) && write_burst_block_ram_wvalid_105)? write_burst_packed_ram_wdata_114 : 'hx;
  assign ram_w8_l4096_id0_1_1_wenable = ((write_burst_packed_fsm_2 == 1) && write_burst_block_ram_wvalid_105)? 1'd1 : 0;
  assign ram_w8_l4096_id0_1_1_enable = ((write_burst_packed_fsm_2 == 1) && write_burst_block_ram_wvalid_105)? 1'd1 : 0;
  wire [10-1:0] write_burst_packed_ram_addr_115;
  assign write_burst_packed_ram_addr_115 = write_burst_packed_addr_107 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_116;
  assign write_burst_packed_ram_wdata_116 = _maxi_rdata_sb_0 >> 16;
  assign ram_w8_l4096_id0_2_1_addr = ((write_burst_packed_fsm_2 == 1) && write_burst_block_ram_wvalid_105)? write_burst_packed_ram_addr_115 : 'hx;
  assign ram_w8_l4096_id0_2_1_wdata = ((write_burst_packed_fsm_2 == 1) && write_burst_block_ram_wvalid_105)? write_burst_packed_ram_wdata_116 : 'hx;
  assign ram_w8_l4096_id0_2_1_wenable = ((write_burst_packed_fsm_2 == 1) && write_burst_block_ram_wvalid_105)? 1'd1 : 0;
  assign ram_w8_l4096_id0_2_1_enable = ((write_burst_packed_fsm_2 == 1) && write_burst_block_ram_wvalid_105)? 1'd1 : 0;
  wire [10-1:0] write_burst_packed_ram_addr_117;
  assign write_burst_packed_ram_addr_117 = write_burst_packed_addr_107 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_118;
  assign write_burst_packed_ram_wdata_118 = _maxi_rdata_sb_0 >> 24;
  assign ram_w8_l4096_id0_3_1_addr = ((write_burst_packed_fsm_2 == 1) && write_burst_block_ram_wvalid_105)? write_burst_packed_ram_addr_117 : 'hx;
  assign ram_w8_l4096_id0_3_1_wdata = ((write_burst_packed_fsm_2 == 1) && write_burst_block_ram_wvalid_105)? write_burst_packed_ram_wdata_118 : 'hx;
  assign ram_w8_l4096_id0_3_1_wenable = ((write_burst_packed_fsm_2 == 1) && write_burst_block_ram_wvalid_105)? 1'd1 : 0;
  assign ram_w8_l4096_id0_3_1_enable = ((write_burst_packed_fsm_2 == 1) && write_burst_block_ram_wvalid_105)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_119;
  wire write_burst_block_ram_wquit_120;
  reg [32-1:0] write_burst_packed_fsm_3;
  localparam write_burst_packed_fsm_3_init = 0;
  reg [12-1:0] write_burst_packed_addr_121;
  reg [12-1:0] write_burst_packed_stride_122;
  reg [33-1:0] write_burst_packed_length_123;
  reg write_burst_packed_done_124;
  wire [10-1:0] write_burst_packed_ram_addr_125;
  assign write_burst_packed_ram_addr_125 = write_burst_packed_addr_121 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_126;
  assign write_burst_packed_ram_wdata_126 = _maxi_rdata_sb_0 >> 0;
  assign ram_w8_l4096_id1_0_1_addr = ((write_burst_packed_fsm_3 == 1) && write_burst_block_ram_wvalid_119)? write_burst_packed_ram_addr_125 : 'hx;
  assign ram_w8_l4096_id1_0_1_wdata = ((write_burst_packed_fsm_3 == 1) && write_burst_block_ram_wvalid_119)? write_burst_packed_ram_wdata_126 : 'hx;
  assign ram_w8_l4096_id1_0_1_wenable = ((write_burst_packed_fsm_3 == 1) && write_burst_block_ram_wvalid_119)? 1'd1 : 0;
  assign ram_w8_l4096_id1_0_1_enable = ((write_burst_packed_fsm_3 == 1) && write_burst_block_ram_wvalid_119)? 1'd1 : 0;
  wire [10-1:0] write_burst_packed_ram_addr_127;
  assign write_burst_packed_ram_addr_127 = write_burst_packed_addr_121 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_128;
  assign write_burst_packed_ram_wdata_128 = _maxi_rdata_sb_0 >> 8;
  assign ram_w8_l4096_id1_1_1_addr = ((write_burst_packed_fsm_3 == 1) && write_burst_block_ram_wvalid_119)? write_burst_packed_ram_addr_127 : 'hx;
  assign ram_w8_l4096_id1_1_1_wdata = ((write_burst_packed_fsm_3 == 1) && write_burst_block_ram_wvalid_119)? write_burst_packed_ram_wdata_128 : 'hx;
  assign ram_w8_l4096_id1_1_1_wenable = ((write_burst_packed_fsm_3 == 1) && write_burst_block_ram_wvalid_119)? 1'd1 : 0;
  assign ram_w8_l4096_id1_1_1_enable = ((write_burst_packed_fsm_3 == 1) && write_burst_block_ram_wvalid_119)? 1'd1 : 0;
  wire [10-1:0] write_burst_packed_ram_addr_129;
  assign write_burst_packed_ram_addr_129 = write_burst_packed_addr_121 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_130;
  assign write_burst_packed_ram_wdata_130 = _maxi_rdata_sb_0 >> 16;
  assign ram_w8_l4096_id1_2_1_addr = ((write_burst_packed_fsm_3 == 1) && write_burst_block_ram_wvalid_119)? write_burst_packed_ram_addr_129 : 'hx;
  assign ram_w8_l4096_id1_2_1_wdata = ((write_burst_packed_fsm_3 == 1) && write_burst_block_ram_wvalid_119)? write_burst_packed_ram_wdata_130 : 'hx;
  assign ram_w8_l4096_id1_2_1_wenable = ((write_burst_packed_fsm_3 == 1) && write_burst_block_ram_wvalid_119)? 1'd1 : 0;
  assign ram_w8_l4096_id1_2_1_enable = ((write_burst_packed_fsm_3 == 1) && write_burst_block_ram_wvalid_119)? 1'd1 : 0;
  wire [10-1:0] write_burst_packed_ram_addr_131;
  assign write_burst_packed_ram_addr_131 = write_burst_packed_addr_121 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_132;
  assign write_burst_packed_ram_wdata_132 = _maxi_rdata_sb_0 >> 24;
  assign ram_w8_l4096_id1_3_1_addr = ((write_burst_packed_fsm_3 == 1) && write_burst_block_ram_wvalid_119)? write_burst_packed_ram_addr_131 : 'hx;
  assign ram_w8_l4096_id1_3_1_wdata = ((write_burst_packed_fsm_3 == 1) && write_burst_block_ram_wvalid_119)? write_burst_packed_ram_wdata_132 : 'hx;
  assign ram_w8_l4096_id1_3_1_wenable = ((write_burst_packed_fsm_3 == 1) && write_burst_block_ram_wvalid_119)? 1'd1 : 0;
  assign ram_w8_l4096_id1_3_1_enable = ((write_burst_packed_fsm_3 == 1) && write_burst_block_ram_wvalid_119)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_133;
  wire write_burst_block_ram_wquit_134;
  reg [32-1:0] write_burst_packed_fsm_4;
  localparam write_burst_packed_fsm_4_init = 0;
  reg [12-1:0] write_burst_packed_addr_135;
  reg [12-1:0] write_burst_packed_stride_136;
  reg [33-1:0] write_burst_packed_length_137;
  reg write_burst_packed_done_138;
  wire [10-1:0] write_burst_packed_ram_addr_139;
  assign write_burst_packed_ram_addr_139 = write_burst_packed_addr_135 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_140;
  assign write_burst_packed_ram_wdata_140 = _maxi_rdata_sb_0 >> 0;
  assign ram_w8_l4096_id2_0_1_addr = ((write_burst_packed_fsm_4 == 1) && write_burst_block_ram_wvalid_133)? write_burst_packed_ram_addr_139 : 'hx;
  assign ram_w8_l4096_id2_0_1_wdata = ((write_burst_packed_fsm_4 == 1) && write_burst_block_ram_wvalid_133)? write_burst_packed_ram_wdata_140 : 'hx;
  assign ram_w8_l4096_id2_0_1_wenable = ((write_burst_packed_fsm_4 == 1) && write_burst_block_ram_wvalid_133)? 1'd1 : 0;
  assign ram_w8_l4096_id2_0_1_enable = ((write_burst_packed_fsm_4 == 1) && write_burst_block_ram_wvalid_133)? 1'd1 : 0;
  wire [10-1:0] write_burst_packed_ram_addr_141;
  assign write_burst_packed_ram_addr_141 = write_burst_packed_addr_135 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_142;
  assign write_burst_packed_ram_wdata_142 = _maxi_rdata_sb_0 >> 8;
  assign ram_w8_l4096_id2_1_1_addr = ((write_burst_packed_fsm_4 == 1) && write_burst_block_ram_wvalid_133)? write_burst_packed_ram_addr_141 : 'hx;
  assign ram_w8_l4096_id2_1_1_wdata = ((write_burst_packed_fsm_4 == 1) && write_burst_block_ram_wvalid_133)? write_burst_packed_ram_wdata_142 : 'hx;
  assign ram_w8_l4096_id2_1_1_wenable = ((write_burst_packed_fsm_4 == 1) && write_burst_block_ram_wvalid_133)? 1'd1 : 0;
  assign ram_w8_l4096_id2_1_1_enable = ((write_burst_packed_fsm_4 == 1) && write_burst_block_ram_wvalid_133)? 1'd1 : 0;
  wire [10-1:0] write_burst_packed_ram_addr_143;
  assign write_burst_packed_ram_addr_143 = write_burst_packed_addr_135 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_144;
  assign write_burst_packed_ram_wdata_144 = _maxi_rdata_sb_0 >> 16;
  assign ram_w8_l4096_id2_2_1_addr = ((write_burst_packed_fsm_4 == 1) && write_burst_block_ram_wvalid_133)? write_burst_packed_ram_addr_143 : 'hx;
  assign ram_w8_l4096_id2_2_1_wdata = ((write_burst_packed_fsm_4 == 1) && write_burst_block_ram_wvalid_133)? write_burst_packed_ram_wdata_144 : 'hx;
  assign ram_w8_l4096_id2_2_1_wenable = ((write_burst_packed_fsm_4 == 1) && write_burst_block_ram_wvalid_133)? 1'd1 : 0;
  assign ram_w8_l4096_id2_2_1_enable = ((write_burst_packed_fsm_4 == 1) && write_burst_block_ram_wvalid_133)? 1'd1 : 0;
  wire [10-1:0] write_burst_packed_ram_addr_145;
  assign write_burst_packed_ram_addr_145 = write_burst_packed_addr_135 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_146;
  assign write_burst_packed_ram_wdata_146 = _maxi_rdata_sb_0 >> 24;
  assign ram_w8_l4096_id2_3_1_addr = ((write_burst_packed_fsm_4 == 1) && write_burst_block_ram_wvalid_133)? write_burst_packed_ram_addr_145 : 'hx;
  assign ram_w8_l4096_id2_3_1_wdata = ((write_burst_packed_fsm_4 == 1) && write_burst_block_ram_wvalid_133)? write_burst_packed_ram_wdata_146 : 'hx;
  assign ram_w8_l4096_id2_3_1_wenable = ((write_burst_packed_fsm_4 == 1) && write_burst_block_ram_wvalid_133)? 1'd1 : 0;
  assign ram_w8_l4096_id2_3_1_enable = ((write_burst_packed_fsm_4 == 1) && write_burst_block_ram_wvalid_133)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_147;
  wire write_burst_block_ram_wquit_148;
  reg [32-1:0] write_burst_packed_fsm_5;
  localparam write_burst_packed_fsm_5_init = 0;
  reg [12-1:0] write_burst_packed_addr_149;
  reg [12-1:0] write_burst_packed_stride_150;
  reg [33-1:0] write_burst_packed_length_151;
  reg write_burst_packed_done_152;
  wire [10-1:0] write_burst_packed_ram_addr_153;
  assign write_burst_packed_ram_addr_153 = write_burst_packed_addr_149 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_154;
  assign write_burst_packed_ram_wdata_154 = _maxi_rdata_sb_0 >> 0;
  assign ram_w8_l4096_id3_0_1_addr = ((write_burst_packed_fsm_5 == 1) && write_burst_block_ram_wvalid_147)? write_burst_packed_ram_addr_153 : 'hx;
  assign ram_w8_l4096_id3_0_1_wdata = ((write_burst_packed_fsm_5 == 1) && write_burst_block_ram_wvalid_147)? write_burst_packed_ram_wdata_154 : 'hx;
  assign ram_w8_l4096_id3_0_1_wenable = ((write_burst_packed_fsm_5 == 1) && write_burst_block_ram_wvalid_147)? 1'd1 : 0;
  assign ram_w8_l4096_id3_0_1_enable = ((write_burst_packed_fsm_5 == 1) && write_burst_block_ram_wvalid_147)? 1'd1 : 0;
  wire [10-1:0] write_burst_packed_ram_addr_155;
  assign write_burst_packed_ram_addr_155 = write_burst_packed_addr_149 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_156;
  assign write_burst_packed_ram_wdata_156 = _maxi_rdata_sb_0 >> 8;
  assign ram_w8_l4096_id3_1_1_addr = ((write_burst_packed_fsm_5 == 1) && write_burst_block_ram_wvalid_147)? write_burst_packed_ram_addr_155 : 'hx;
  assign ram_w8_l4096_id3_1_1_wdata = ((write_burst_packed_fsm_5 == 1) && write_burst_block_ram_wvalid_147)? write_burst_packed_ram_wdata_156 : 'hx;
  assign ram_w8_l4096_id3_1_1_wenable = ((write_burst_packed_fsm_5 == 1) && write_burst_block_ram_wvalid_147)? 1'd1 : 0;
  assign ram_w8_l4096_id3_1_1_enable = ((write_burst_packed_fsm_5 == 1) && write_burst_block_ram_wvalid_147)? 1'd1 : 0;
  wire [10-1:0] write_burst_packed_ram_addr_157;
  assign write_burst_packed_ram_addr_157 = write_burst_packed_addr_149 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_158;
  assign write_burst_packed_ram_wdata_158 = _maxi_rdata_sb_0 >> 16;
  assign ram_w8_l4096_id3_2_1_addr = ((write_burst_packed_fsm_5 == 1) && write_burst_block_ram_wvalid_147)? write_burst_packed_ram_addr_157 : 'hx;
  assign ram_w8_l4096_id3_2_1_wdata = ((write_burst_packed_fsm_5 == 1) && write_burst_block_ram_wvalid_147)? write_burst_packed_ram_wdata_158 : 'hx;
  assign ram_w8_l4096_id3_2_1_wenable = ((write_burst_packed_fsm_5 == 1) && write_burst_block_ram_wvalid_147)? 1'd1 : 0;
  assign ram_w8_l4096_id3_2_1_enable = ((write_burst_packed_fsm_5 == 1) && write_burst_block_ram_wvalid_147)? 1'd1 : 0;
  wire [10-1:0] write_burst_packed_ram_addr_159;
  assign write_burst_packed_ram_addr_159 = write_burst_packed_addr_149 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_160;
  assign write_burst_packed_ram_wdata_160 = _maxi_rdata_sb_0 >> 24;
  assign ram_w8_l4096_id3_3_1_addr = ((write_burst_packed_fsm_5 == 1) && write_burst_block_ram_wvalid_147)? write_burst_packed_ram_addr_159 : 'hx;
  assign ram_w8_l4096_id3_3_1_wdata = ((write_burst_packed_fsm_5 == 1) && write_burst_block_ram_wvalid_147)? write_burst_packed_ram_wdata_160 : 'hx;
  assign ram_w8_l4096_id3_3_1_wenable = ((write_burst_packed_fsm_5 == 1) && write_burst_block_ram_wvalid_147)? 1'd1 : 0;
  assign ram_w8_l4096_id3_3_1_enable = ((write_burst_packed_fsm_5 == 1) && write_burst_block_ram_wvalid_147)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_161;
  wire write_burst_block_ram_wquit_162;
  reg [32-1:0] write_burst_packed_fsm_6;
  localparam write_burst_packed_fsm_6_init = 0;
  reg [12-1:0] write_burst_packed_addr_163;
  reg [12-1:0] write_burst_packed_stride_164;
  reg [33-1:0] write_burst_packed_length_165;
  reg write_burst_packed_done_166;
  wire [10-1:0] write_burst_packed_ram_addr_167;
  assign write_burst_packed_ram_addr_167 = write_burst_packed_addr_163 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_168;
  assign write_burst_packed_ram_wdata_168 = _maxi_rdata_sb_0 >> 0;
  assign ram_w8_l4096_id4_0_1_addr = ((write_burst_packed_fsm_6 == 1) && write_burst_block_ram_wvalid_161)? write_burst_packed_ram_addr_167 : 'hx;
  assign ram_w8_l4096_id4_0_1_wdata = ((write_burst_packed_fsm_6 == 1) && write_burst_block_ram_wvalid_161)? write_burst_packed_ram_wdata_168 : 'hx;
  assign ram_w8_l4096_id4_0_1_wenable = ((write_burst_packed_fsm_6 == 1) && write_burst_block_ram_wvalid_161)? 1'd1 : 0;
  assign ram_w8_l4096_id4_0_1_enable = ((write_burst_packed_fsm_6 == 1) && write_burst_block_ram_wvalid_161)? 1'd1 : 0;
  wire [10-1:0] write_burst_packed_ram_addr_169;
  assign write_burst_packed_ram_addr_169 = write_burst_packed_addr_163 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_170;
  assign write_burst_packed_ram_wdata_170 = _maxi_rdata_sb_0 >> 8;
  assign ram_w8_l4096_id4_1_1_addr = ((write_burst_packed_fsm_6 == 1) && write_burst_block_ram_wvalid_161)? write_burst_packed_ram_addr_169 : 'hx;
  assign ram_w8_l4096_id4_1_1_wdata = ((write_burst_packed_fsm_6 == 1) && write_burst_block_ram_wvalid_161)? write_burst_packed_ram_wdata_170 : 'hx;
  assign ram_w8_l4096_id4_1_1_wenable = ((write_burst_packed_fsm_6 == 1) && write_burst_block_ram_wvalid_161)? 1'd1 : 0;
  assign ram_w8_l4096_id4_1_1_enable = ((write_burst_packed_fsm_6 == 1) && write_burst_block_ram_wvalid_161)? 1'd1 : 0;
  wire [10-1:0] write_burst_packed_ram_addr_171;
  assign write_burst_packed_ram_addr_171 = write_burst_packed_addr_163 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_172;
  assign write_burst_packed_ram_wdata_172 = _maxi_rdata_sb_0 >> 16;
  assign ram_w8_l4096_id4_2_1_addr = ((write_burst_packed_fsm_6 == 1) && write_burst_block_ram_wvalid_161)? write_burst_packed_ram_addr_171 : 'hx;
  assign ram_w8_l4096_id4_2_1_wdata = ((write_burst_packed_fsm_6 == 1) && write_burst_block_ram_wvalid_161)? write_burst_packed_ram_wdata_172 : 'hx;
  assign ram_w8_l4096_id4_2_1_wenable = ((write_burst_packed_fsm_6 == 1) && write_burst_block_ram_wvalid_161)? 1'd1 : 0;
  assign ram_w8_l4096_id4_2_1_enable = ((write_burst_packed_fsm_6 == 1) && write_burst_block_ram_wvalid_161)? 1'd1 : 0;
  wire [10-1:0] write_burst_packed_ram_addr_173;
  assign write_burst_packed_ram_addr_173 = write_burst_packed_addr_163 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_174;
  assign write_burst_packed_ram_wdata_174 = _maxi_rdata_sb_0 >> 24;
  assign ram_w8_l4096_id4_3_1_addr = ((write_burst_packed_fsm_6 == 1) && write_burst_block_ram_wvalid_161)? write_burst_packed_ram_addr_173 : 'hx;
  assign ram_w8_l4096_id4_3_1_wdata = ((write_burst_packed_fsm_6 == 1) && write_burst_block_ram_wvalid_161)? write_burst_packed_ram_wdata_174 : 'hx;
  assign ram_w8_l4096_id4_3_1_wenable = ((write_burst_packed_fsm_6 == 1) && write_burst_block_ram_wvalid_161)? 1'd1 : 0;
  assign ram_w8_l4096_id4_3_1_enable = ((write_burst_packed_fsm_6 == 1) && write_burst_block_ram_wvalid_161)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_175;
  wire write_burst_block_ram_wquit_176;
  reg [32-1:0] write_burst_packed_fsm_7;
  localparam write_burst_packed_fsm_7_init = 0;
  reg [12-1:0] write_burst_packed_addr_177;
  reg [12-1:0] write_burst_packed_stride_178;
  reg [33-1:0] write_burst_packed_length_179;
  reg write_burst_packed_done_180;
  wire [10-1:0] write_burst_packed_ram_addr_181;
  assign write_burst_packed_ram_addr_181 = write_burst_packed_addr_177 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_182;
  assign write_burst_packed_ram_wdata_182 = _maxi_rdata_sb_0 >> 0;
  assign ram_w8_l4096_id5_0_1_addr = ((write_burst_packed_fsm_7 == 1) && write_burst_block_ram_wvalid_175)? write_burst_packed_ram_addr_181 : 'hx;
  assign ram_w8_l4096_id5_0_1_wdata = ((write_burst_packed_fsm_7 == 1) && write_burst_block_ram_wvalid_175)? write_burst_packed_ram_wdata_182 : 'hx;
  assign ram_w8_l4096_id5_0_1_wenable = ((write_burst_packed_fsm_7 == 1) && write_burst_block_ram_wvalid_175)? 1'd1 : 0;
  assign ram_w8_l4096_id5_0_1_enable = ((write_burst_packed_fsm_7 == 1) && write_burst_block_ram_wvalid_175)? 1'd1 : 0;
  wire [10-1:0] write_burst_packed_ram_addr_183;
  assign write_burst_packed_ram_addr_183 = write_burst_packed_addr_177 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_184;
  assign write_burst_packed_ram_wdata_184 = _maxi_rdata_sb_0 >> 8;
  assign ram_w8_l4096_id5_1_1_addr = ((write_burst_packed_fsm_7 == 1) && write_burst_block_ram_wvalid_175)? write_burst_packed_ram_addr_183 : 'hx;
  assign ram_w8_l4096_id5_1_1_wdata = ((write_burst_packed_fsm_7 == 1) && write_burst_block_ram_wvalid_175)? write_burst_packed_ram_wdata_184 : 'hx;
  assign ram_w8_l4096_id5_1_1_wenable = ((write_burst_packed_fsm_7 == 1) && write_burst_block_ram_wvalid_175)? 1'd1 : 0;
  assign ram_w8_l4096_id5_1_1_enable = ((write_burst_packed_fsm_7 == 1) && write_burst_block_ram_wvalid_175)? 1'd1 : 0;
  wire [10-1:0] write_burst_packed_ram_addr_185;
  assign write_burst_packed_ram_addr_185 = write_burst_packed_addr_177 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_186;
  assign write_burst_packed_ram_wdata_186 = _maxi_rdata_sb_0 >> 16;
  assign ram_w8_l4096_id5_2_1_addr = ((write_burst_packed_fsm_7 == 1) && write_burst_block_ram_wvalid_175)? write_burst_packed_ram_addr_185 : 'hx;
  assign ram_w8_l4096_id5_2_1_wdata = ((write_burst_packed_fsm_7 == 1) && write_burst_block_ram_wvalid_175)? write_burst_packed_ram_wdata_186 : 'hx;
  assign ram_w8_l4096_id5_2_1_wenable = ((write_burst_packed_fsm_7 == 1) && write_burst_block_ram_wvalid_175)? 1'd1 : 0;
  assign ram_w8_l4096_id5_2_1_enable = ((write_burst_packed_fsm_7 == 1) && write_burst_block_ram_wvalid_175)? 1'd1 : 0;
  wire [10-1:0] write_burst_packed_ram_addr_187;
  assign write_burst_packed_ram_addr_187 = write_burst_packed_addr_177 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_188;
  assign write_burst_packed_ram_wdata_188 = _maxi_rdata_sb_0 >> 24;
  assign ram_w8_l4096_id5_3_1_addr = ((write_burst_packed_fsm_7 == 1) && write_burst_block_ram_wvalid_175)? write_burst_packed_ram_addr_187 : 'hx;
  assign ram_w8_l4096_id5_3_1_wdata = ((write_burst_packed_fsm_7 == 1) && write_burst_block_ram_wvalid_175)? write_burst_packed_ram_wdata_188 : 'hx;
  assign ram_w8_l4096_id5_3_1_wenable = ((write_burst_packed_fsm_7 == 1) && write_burst_block_ram_wvalid_175)? 1'd1 : 0;
  assign ram_w8_l4096_id5_3_1_enable = ((write_burst_packed_fsm_7 == 1) && write_burst_block_ram_wvalid_175)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_189;
  wire write_burst_block_ram_wquit_190;
  reg [32-1:0] write_burst_packed_fsm_8;
  localparam write_burst_packed_fsm_8_init = 0;
  reg [12-1:0] write_burst_packed_addr_191;
  reg [12-1:0] write_burst_packed_stride_192;
  reg [33-1:0] write_burst_packed_length_193;
  reg write_burst_packed_done_194;
  wire [10-1:0] write_burst_packed_ram_addr_195;
  assign write_burst_packed_ram_addr_195 = write_burst_packed_addr_191 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_196;
  assign write_burst_packed_ram_wdata_196 = _maxi_rdata_sb_0 >> 0;
  assign ram_w8_l4096_id6_0_1_addr = ((write_burst_packed_fsm_8 == 1) && write_burst_block_ram_wvalid_189)? write_burst_packed_ram_addr_195 : 'hx;
  assign ram_w8_l4096_id6_0_1_wdata = ((write_burst_packed_fsm_8 == 1) && write_burst_block_ram_wvalid_189)? write_burst_packed_ram_wdata_196 : 'hx;
  assign ram_w8_l4096_id6_0_1_wenable = ((write_burst_packed_fsm_8 == 1) && write_burst_block_ram_wvalid_189)? 1'd1 : 0;
  assign ram_w8_l4096_id6_0_1_enable = ((write_burst_packed_fsm_8 == 1) && write_burst_block_ram_wvalid_189)? 1'd1 : 0;
  wire [10-1:0] write_burst_packed_ram_addr_197;
  assign write_burst_packed_ram_addr_197 = write_burst_packed_addr_191 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_198;
  assign write_burst_packed_ram_wdata_198 = _maxi_rdata_sb_0 >> 8;
  assign ram_w8_l4096_id6_1_1_addr = ((write_burst_packed_fsm_8 == 1) && write_burst_block_ram_wvalid_189)? write_burst_packed_ram_addr_197 : 'hx;
  assign ram_w8_l4096_id6_1_1_wdata = ((write_burst_packed_fsm_8 == 1) && write_burst_block_ram_wvalid_189)? write_burst_packed_ram_wdata_198 : 'hx;
  assign ram_w8_l4096_id6_1_1_wenable = ((write_burst_packed_fsm_8 == 1) && write_burst_block_ram_wvalid_189)? 1'd1 : 0;
  assign ram_w8_l4096_id6_1_1_enable = ((write_burst_packed_fsm_8 == 1) && write_burst_block_ram_wvalid_189)? 1'd1 : 0;
  wire [10-1:0] write_burst_packed_ram_addr_199;
  assign write_burst_packed_ram_addr_199 = write_burst_packed_addr_191 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_200;
  assign write_burst_packed_ram_wdata_200 = _maxi_rdata_sb_0 >> 16;
  assign ram_w8_l4096_id6_2_1_addr = ((write_burst_packed_fsm_8 == 1) && write_burst_block_ram_wvalid_189)? write_burst_packed_ram_addr_199 : 'hx;
  assign ram_w8_l4096_id6_2_1_wdata = ((write_burst_packed_fsm_8 == 1) && write_burst_block_ram_wvalid_189)? write_burst_packed_ram_wdata_200 : 'hx;
  assign ram_w8_l4096_id6_2_1_wenable = ((write_burst_packed_fsm_8 == 1) && write_burst_block_ram_wvalid_189)? 1'd1 : 0;
  assign ram_w8_l4096_id6_2_1_enable = ((write_burst_packed_fsm_8 == 1) && write_burst_block_ram_wvalid_189)? 1'd1 : 0;
  wire [10-1:0] write_burst_packed_ram_addr_201;
  assign write_burst_packed_ram_addr_201 = write_burst_packed_addr_191 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_202;
  assign write_burst_packed_ram_wdata_202 = _maxi_rdata_sb_0 >> 24;
  assign ram_w8_l4096_id6_3_1_addr = ((write_burst_packed_fsm_8 == 1) && write_burst_block_ram_wvalid_189)? write_burst_packed_ram_addr_201 : 'hx;
  assign ram_w8_l4096_id6_3_1_wdata = ((write_burst_packed_fsm_8 == 1) && write_burst_block_ram_wvalid_189)? write_burst_packed_ram_wdata_202 : 'hx;
  assign ram_w8_l4096_id6_3_1_wenable = ((write_burst_packed_fsm_8 == 1) && write_burst_block_ram_wvalid_189)? 1'd1 : 0;
  assign ram_w8_l4096_id6_3_1_enable = ((write_burst_packed_fsm_8 == 1) && write_burst_block_ram_wvalid_189)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_203;
  wire write_burst_block_ram_wquit_204;
  reg [32-1:0] write_burst_packed_fsm_9;
  localparam write_burst_packed_fsm_9_init = 0;
  reg [12-1:0] write_burst_packed_addr_205;
  reg [12-1:0] write_burst_packed_stride_206;
  reg [33-1:0] write_burst_packed_length_207;
  reg write_burst_packed_done_208;
  wire [10-1:0] write_burst_packed_ram_addr_209;
  assign write_burst_packed_ram_addr_209 = write_burst_packed_addr_205 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_210;
  assign write_burst_packed_ram_wdata_210 = _maxi_rdata_sb_0 >> 0;
  assign ram_w8_l4096_id7_0_1_addr = ((write_burst_packed_fsm_9 == 1) && write_burst_block_ram_wvalid_203)? write_burst_packed_ram_addr_209 : 'hx;
  assign ram_w8_l4096_id7_0_1_wdata = ((write_burst_packed_fsm_9 == 1) && write_burst_block_ram_wvalid_203)? write_burst_packed_ram_wdata_210 : 'hx;
  assign ram_w8_l4096_id7_0_1_wenable = ((write_burst_packed_fsm_9 == 1) && write_burst_block_ram_wvalid_203)? 1'd1 : 0;
  assign ram_w8_l4096_id7_0_1_enable = ((write_burst_packed_fsm_9 == 1) && write_burst_block_ram_wvalid_203)? 1'd1 : 0;
  wire [10-1:0] write_burst_packed_ram_addr_211;
  assign write_burst_packed_ram_addr_211 = write_burst_packed_addr_205 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_212;
  assign write_burst_packed_ram_wdata_212 = _maxi_rdata_sb_0 >> 8;
  assign ram_w8_l4096_id7_1_1_addr = ((write_burst_packed_fsm_9 == 1) && write_burst_block_ram_wvalid_203)? write_burst_packed_ram_addr_211 : 'hx;
  assign ram_w8_l4096_id7_1_1_wdata = ((write_burst_packed_fsm_9 == 1) && write_burst_block_ram_wvalid_203)? write_burst_packed_ram_wdata_212 : 'hx;
  assign ram_w8_l4096_id7_1_1_wenable = ((write_burst_packed_fsm_9 == 1) && write_burst_block_ram_wvalid_203)? 1'd1 : 0;
  assign ram_w8_l4096_id7_1_1_enable = ((write_burst_packed_fsm_9 == 1) && write_burst_block_ram_wvalid_203)? 1'd1 : 0;
  wire [10-1:0] write_burst_packed_ram_addr_213;
  assign write_burst_packed_ram_addr_213 = write_burst_packed_addr_205 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_214;
  assign write_burst_packed_ram_wdata_214 = _maxi_rdata_sb_0 >> 16;
  assign ram_w8_l4096_id7_2_1_addr = ((write_burst_packed_fsm_9 == 1) && write_burst_block_ram_wvalid_203)? write_burst_packed_ram_addr_213 : 'hx;
  assign ram_w8_l4096_id7_2_1_wdata = ((write_burst_packed_fsm_9 == 1) && write_burst_block_ram_wvalid_203)? write_burst_packed_ram_wdata_214 : 'hx;
  assign ram_w8_l4096_id7_2_1_wenable = ((write_burst_packed_fsm_9 == 1) && write_burst_block_ram_wvalid_203)? 1'd1 : 0;
  assign ram_w8_l4096_id7_2_1_enable = ((write_burst_packed_fsm_9 == 1) && write_burst_block_ram_wvalid_203)? 1'd1 : 0;
  wire [10-1:0] write_burst_packed_ram_addr_215;
  assign write_burst_packed_ram_addr_215 = write_burst_packed_addr_205 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_216;
  assign write_burst_packed_ram_wdata_216 = _maxi_rdata_sb_0 >> 24;
  assign ram_w8_l4096_id7_3_1_addr = ((write_burst_packed_fsm_9 == 1) && write_burst_block_ram_wvalid_203)? write_burst_packed_ram_addr_215 : 'hx;
  assign ram_w8_l4096_id7_3_1_wdata = ((write_burst_packed_fsm_9 == 1) && write_burst_block_ram_wvalid_203)? write_burst_packed_ram_wdata_216 : 'hx;
  assign ram_w8_l4096_id7_3_1_wenable = ((write_burst_packed_fsm_9 == 1) && write_burst_block_ram_wvalid_203)? 1'd1 : 0;
  assign ram_w8_l4096_id7_3_1_enable = ((write_burst_packed_fsm_9 == 1) && write_burst_block_ram_wvalid_203)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_217;
  wire write_burst_block_ram_wquit_218;
  reg [32-1:0] write_burst_packed_fsm_10;
  localparam write_burst_packed_fsm_10_init = 0;
  reg [12-1:0] write_burst_packed_addr_219;
  reg [12-1:0] write_burst_packed_stride_220;
  reg [33-1:0] write_burst_packed_length_221;
  reg write_burst_packed_done_222;
  wire [10-1:0] write_burst_packed_ram_addr_223;
  assign write_burst_packed_ram_addr_223 = write_burst_packed_addr_219 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_224;
  assign write_burst_packed_ram_wdata_224 = _maxi_rdata_sb_0 >> 0;
  assign ram_w8_l4096_id8_0_1_addr = ((write_burst_packed_fsm_10 == 1) && write_burst_block_ram_wvalid_217)? write_burst_packed_ram_addr_223 : 'hx;
  assign ram_w8_l4096_id8_0_1_wdata = ((write_burst_packed_fsm_10 == 1) && write_burst_block_ram_wvalid_217)? write_burst_packed_ram_wdata_224 : 'hx;
  assign ram_w8_l4096_id8_0_1_wenable = ((write_burst_packed_fsm_10 == 1) && write_burst_block_ram_wvalid_217)? 1'd1 : 0;
  assign ram_w8_l4096_id8_0_1_enable = ((write_burst_packed_fsm_10 == 1) && write_burst_block_ram_wvalid_217)? 1'd1 : 0;
  wire [10-1:0] write_burst_packed_ram_addr_225;
  assign write_burst_packed_ram_addr_225 = write_burst_packed_addr_219 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_226;
  assign write_burst_packed_ram_wdata_226 = _maxi_rdata_sb_0 >> 8;
  assign ram_w8_l4096_id8_1_1_addr = ((write_burst_packed_fsm_10 == 1) && write_burst_block_ram_wvalid_217)? write_burst_packed_ram_addr_225 : 'hx;
  assign ram_w8_l4096_id8_1_1_wdata = ((write_burst_packed_fsm_10 == 1) && write_burst_block_ram_wvalid_217)? write_burst_packed_ram_wdata_226 : 'hx;
  assign ram_w8_l4096_id8_1_1_wenable = ((write_burst_packed_fsm_10 == 1) && write_burst_block_ram_wvalid_217)? 1'd1 : 0;
  assign ram_w8_l4096_id8_1_1_enable = ((write_burst_packed_fsm_10 == 1) && write_burst_block_ram_wvalid_217)? 1'd1 : 0;
  wire [10-1:0] write_burst_packed_ram_addr_227;
  assign write_burst_packed_ram_addr_227 = write_burst_packed_addr_219 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_228;
  assign write_burst_packed_ram_wdata_228 = _maxi_rdata_sb_0 >> 16;
  assign ram_w8_l4096_id8_2_1_addr = ((write_burst_packed_fsm_10 == 1) && write_burst_block_ram_wvalid_217)? write_burst_packed_ram_addr_227 : 'hx;
  assign ram_w8_l4096_id8_2_1_wdata = ((write_burst_packed_fsm_10 == 1) && write_burst_block_ram_wvalid_217)? write_burst_packed_ram_wdata_228 : 'hx;
  assign ram_w8_l4096_id8_2_1_wenable = ((write_burst_packed_fsm_10 == 1) && write_burst_block_ram_wvalid_217)? 1'd1 : 0;
  assign ram_w8_l4096_id8_2_1_enable = ((write_burst_packed_fsm_10 == 1) && write_burst_block_ram_wvalid_217)? 1'd1 : 0;
  wire [10-1:0] write_burst_packed_ram_addr_229;
  assign write_burst_packed_ram_addr_229 = write_burst_packed_addr_219 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_230;
  assign write_burst_packed_ram_wdata_230 = _maxi_rdata_sb_0 >> 24;
  assign ram_w8_l4096_id8_3_1_addr = ((write_burst_packed_fsm_10 == 1) && write_burst_block_ram_wvalid_217)? write_burst_packed_ram_addr_229 : 'hx;
  assign ram_w8_l4096_id8_3_1_wdata = ((write_burst_packed_fsm_10 == 1) && write_burst_block_ram_wvalid_217)? write_burst_packed_ram_wdata_230 : 'hx;
  assign ram_w8_l4096_id8_3_1_wenable = ((write_burst_packed_fsm_10 == 1) && write_burst_block_ram_wvalid_217)? 1'd1 : 0;
  assign ram_w8_l4096_id8_3_1_enable = ((write_burst_packed_fsm_10 == 1) && write_burst_block_ram_wvalid_217)? 1'd1 : 0;
  reg [32-1:0] write_burst_block_fsm_11;
  localparam write_burst_block_fsm_11_init = 0;
  reg [33-1:0] write_burst_block_length_231;
  reg [32-1:0] write_burst_block_blocksize_232;
  reg write_burst_block_done_233;
  reg [32-1:0] write_burst_block_count_234;
  assign write_burst_block_ram_wvalid_105 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_11 == 1);
  assign write_burst_block_ram_wquit_106 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_231 <= 1);
  assign write_burst_block_ram_wvalid_119 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_11 == 2);
  assign write_burst_block_ram_wquit_120 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_231 <= 1);
  assign write_burst_block_ram_wvalid_133 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_11 == 3);
  assign write_burst_block_ram_wquit_134 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_231 <= 1);
  assign write_burst_block_ram_wvalid_147 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_11 == 4);
  assign write_burst_block_ram_wquit_148 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_231 <= 1);
  assign write_burst_block_ram_wvalid_161 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_11 == 5);
  assign write_burst_block_ram_wquit_162 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_231 <= 1);
  assign write_burst_block_ram_wvalid_175 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_11 == 6);
  assign write_burst_block_ram_wquit_176 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_231 <= 1);
  assign write_burst_block_ram_wvalid_189 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_11 == 7);
  assign write_burst_block_ram_wquit_190 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_231 <= 1);
  assign write_burst_block_ram_wvalid_203 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_11 == 8);
  assign write_burst_block_ram_wquit_204 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_231 <= 1);
  assign write_burst_block_ram_wvalid_217 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_11 == 9);
  assign write_burst_block_ram_wquit_218 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_231 <= 1);
  wire [32-1:0] conv2d_24_mux_act_gaddr_0;
  assign conv2d_24_mux_act_gaddr_0 = (conv2d_24_row_select == 0)? conv2d_24_arg_objaddr_0 + (conv2d_24_act_base_offset + cparam_conv2d_24_act_offset_values_0) : 
                                     (conv2d_24_row_select == 1)? conv2d_24_arg_objaddr_0 + (conv2d_24_act_base_offset + cparam_conv2d_24_act_offset_values_2) : 
                                     (conv2d_24_row_select == 2)? conv2d_24_arg_objaddr_0 + (conv2d_24_act_base_offset + cparam_conv2d_24_act_offset_values_1) : 1'd0;
  wire [32-1:0] conv2d_24_mux_act_gaddr_1;
  assign conv2d_24_mux_act_gaddr_1 = (conv2d_24_row_select == 0)? conv2d_24_arg_objaddr_0 + (conv2d_24_act_base_offset + cparam_conv2d_24_act_offset_values_1) : 
                                     (conv2d_24_row_select == 1)? conv2d_24_arg_objaddr_0 + (conv2d_24_act_base_offset + cparam_conv2d_24_act_offset_values_0) : 
                                     (conv2d_24_row_select == 2)? conv2d_24_arg_objaddr_0 + (conv2d_24_act_base_offset + cparam_conv2d_24_act_offset_values_2) : 1'd0;
  wire [32-1:0] conv2d_24_mux_act_gaddr_2;
  assign conv2d_24_mux_act_gaddr_2 = (conv2d_24_row_select == 0)? conv2d_24_arg_objaddr_0 + (conv2d_24_act_base_offset + cparam_conv2d_24_act_offset_values_2) : 
                                     (conv2d_24_row_select == 1)? conv2d_24_arg_objaddr_0 + (conv2d_24_act_base_offset + cparam_conv2d_24_act_offset_values_1) : 
                                     (conv2d_24_row_select == 2)? conv2d_24_arg_objaddr_0 + (conv2d_24_act_base_offset + cparam_conv2d_24_act_offset_values_0) : 1'd0;
  wire conv2d_24_dma_pad_mask_0;
  assign conv2d_24_dma_pad_mask_0 = (conv2d_24_row_count + 0 < cparam_conv2d_24_pad_row_top) || (conv2d_24_row_count + 0 >= cparam_conv2d_24_act_num_row + cparam_conv2d_24_pad_row_top);
  wire conv2d_24_dma_pad_mask_1;
  assign conv2d_24_dma_pad_mask_1 = (conv2d_24_row_count + 1 < cparam_conv2d_24_pad_row_top) || (conv2d_24_row_count + 1 >= cparam_conv2d_24_act_num_row + cparam_conv2d_24_pad_row_top);
  wire conv2d_24_dma_pad_mask_2;
  assign conv2d_24_dma_pad_mask_2 = (conv2d_24_row_count + 2 < cparam_conv2d_24_pad_row_top) || (conv2d_24_row_count + 2 >= cparam_conv2d_24_act_num_row + cparam_conv2d_24_pad_row_top);
  wire conv2d_24_mux_dma_pad_mask_0;
  assign conv2d_24_mux_dma_pad_mask_0 = (conv2d_24_row_select == 0)? conv2d_24_dma_pad_mask_0 : 
                                        (conv2d_24_row_select == 1)? conv2d_24_dma_pad_mask_2 : 
                                        (conv2d_24_row_select == 2)? conv2d_24_dma_pad_mask_1 : 1'd0;
  wire conv2d_24_mux_dma_pad_mask_1;
  assign conv2d_24_mux_dma_pad_mask_1 = (conv2d_24_row_select == 0)? conv2d_24_dma_pad_mask_1 : 
                                        (conv2d_24_row_select == 1)? conv2d_24_dma_pad_mask_0 : 
                                        (conv2d_24_row_select == 2)? conv2d_24_dma_pad_mask_2 : 1'd0;
  wire conv2d_24_mux_dma_pad_mask_2;
  assign conv2d_24_mux_dma_pad_mask_2 = (conv2d_24_row_select == 0)? conv2d_24_dma_pad_mask_2 : 
                                        (conv2d_24_row_select == 1)? conv2d_24_dma_pad_mask_1 : 
                                        (conv2d_24_row_select == 2)? conv2d_24_dma_pad_mask_0 : 1'd0;
  wire conv2d_24_mux_dma_flag_0;
  assign conv2d_24_mux_dma_flag_0 = (conv2d_24_prev_row_select == 0)? conv2d_24_dma_flag_0 : 
                                    (conv2d_24_prev_row_select == 1)? conv2d_24_dma_flag_2 : 
                                    (conv2d_24_prev_row_select == 2)? conv2d_24_dma_flag_1 : 1'd0;
  wire conv2d_24_mux_dma_flag_1;
  assign conv2d_24_mux_dma_flag_1 = (conv2d_24_prev_row_select == 0)? conv2d_24_dma_flag_1 : 
                                    (conv2d_24_prev_row_select == 1)? conv2d_24_dma_flag_0 : 
                                    (conv2d_24_prev_row_select == 2)? conv2d_24_dma_flag_2 : 1'd0;
  wire conv2d_24_mux_dma_flag_2;
  assign conv2d_24_mux_dma_flag_2 = (conv2d_24_prev_row_select == 0)? conv2d_24_dma_flag_2 : 
                                    (conv2d_24_prev_row_select == 1)? conv2d_24_dma_flag_1 : 
                                    (conv2d_24_prev_row_select == 2)? conv2d_24_dma_flag_0 : 1'd0;
  wire [14-1:0] _dma_write_block_high_local_size_235;
  assign _dma_write_block_high_local_size_235 = cparam_conv2d_24_act_read_size >> 2;
  wire [2-1:0] _dma_write_block_low_local_size_236;
  assign _dma_write_block_low_local_size_236 = cparam_conv2d_24_act_read_size & { 2{ 1'd1 } };
  wire [14-1:0] _dma_write_block_local_size_237;
  assign _dma_write_block_local_size_237 = (_dma_write_block_low_local_size_236 > 0)? _dma_write_block_high_local_size_235 + 1 : _dma_write_block_high_local_size_235;
  wire [10-1:0] _dma_read_block_high_local_blocksize_238;
  assign _dma_read_block_high_local_blocksize_238 = cparam_conv2d_24_act_read_block >> 2;
  wire [3-1:0] _dma_read_block_low_local_blocksize_239;
  assign _dma_read_block_low_local_blocksize_239 = cparam_conv2d_24_act_read_block & { 2{ 1'd1 } };
  wire [10-1:0] _dma_read_block_local_blocksize_240;
  assign _dma_read_block_local_blocksize_240 = (_dma_read_block_low_local_blocksize_239 > 0)? _dma_read_block_high_local_blocksize_238 + 1 : _dma_read_block_high_local_blocksize_238;
  wire [32-1:0] mask_addr_shifted_241;
  assign mask_addr_shifted_241 = conv2d_24_mux_act_gaddr_0 + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_242;
  assign mask_addr_masked_242 = mask_addr_shifted_241 << 2;
  wire write_burst_block_ram_wvalid_243;
  wire write_burst_block_ram_wquit_244;
  reg [32-1:0] write_burst_packed_fsm_12;
  localparam write_burst_packed_fsm_12_init = 0;
  reg [14-1:0] write_burst_packed_addr_245;
  reg [14-1:0] write_burst_packed_stride_246;
  reg [33-1:0] write_burst_packed_length_247;
  reg write_burst_packed_done_248;
  wire [12-1:0] write_burst_packed_ram_addr_249;
  assign write_burst_packed_ram_addr_249 = write_burst_packed_addr_245 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_250;
  assign write_burst_packed_ram_wdata_250 = _maxi_rdata_sb_0 >> 0;
  wire [12-1:0] write_burst_packed_ram_addr_251;
  assign write_burst_packed_ram_addr_251 = write_burst_packed_addr_245 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_252;
  assign write_burst_packed_ram_wdata_252 = _maxi_rdata_sb_0 >> 8;
  wire [12-1:0] write_burst_packed_ram_addr_253;
  assign write_burst_packed_ram_addr_253 = write_burst_packed_addr_245 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_254;
  assign write_burst_packed_ram_wdata_254 = _maxi_rdata_sb_0 >> 16;
  wire [12-1:0] write_burst_packed_ram_addr_255;
  assign write_burst_packed_ram_addr_255 = write_burst_packed_addr_245 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_256;
  assign write_burst_packed_ram_wdata_256 = _maxi_rdata_sb_0 >> 24;
  wire write_burst_block_ram_wvalid_257;
  wire write_burst_block_ram_wquit_258;
  reg [32-1:0] write_burst_packed_fsm_13;
  localparam write_burst_packed_fsm_13_init = 0;
  reg [14-1:0] write_burst_packed_addr_259;
  reg [14-1:0] write_burst_packed_stride_260;
  reg [33-1:0] write_burst_packed_length_261;
  reg write_burst_packed_done_262;
  wire [12-1:0] write_burst_packed_ram_addr_263;
  assign write_burst_packed_ram_addr_263 = write_burst_packed_addr_259 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_264;
  assign write_burst_packed_ram_wdata_264 = _maxi_rdata_sb_0 >> 0;
  assign ram_w8_l16384_id1_0_1_wdata = ((write_burst_packed_fsm_13 == 1) && write_burst_block_ram_wvalid_257)? write_burst_packed_ram_wdata_264 : 'hx;
  assign ram_w8_l16384_id1_0_1_wenable = ((write_burst_packed_fsm_13 == 1) && write_burst_block_ram_wvalid_257)? 1'd1 : 0;
  wire [12-1:0] write_burst_packed_ram_addr_265;
  assign write_burst_packed_ram_addr_265 = write_burst_packed_addr_259 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_266;
  assign write_burst_packed_ram_wdata_266 = _maxi_rdata_sb_0 >> 8;
  assign ram_w8_l16384_id1_1_1_wdata = ((write_burst_packed_fsm_13 == 1) && write_burst_block_ram_wvalid_257)? write_burst_packed_ram_wdata_266 : 'hx;
  assign ram_w8_l16384_id1_1_1_wenable = ((write_burst_packed_fsm_13 == 1) && write_burst_block_ram_wvalid_257)? 1'd1 : 0;
  wire [12-1:0] write_burst_packed_ram_addr_267;
  assign write_burst_packed_ram_addr_267 = write_burst_packed_addr_259 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_268;
  assign write_burst_packed_ram_wdata_268 = _maxi_rdata_sb_0 >> 16;
  assign ram_w8_l16384_id1_2_1_wdata = ((write_burst_packed_fsm_13 == 1) && write_burst_block_ram_wvalid_257)? write_burst_packed_ram_wdata_268 : 'hx;
  assign ram_w8_l16384_id1_2_1_wenable = ((write_burst_packed_fsm_13 == 1) && write_burst_block_ram_wvalid_257)? 1'd1 : 0;
  wire [12-1:0] write_burst_packed_ram_addr_269;
  assign write_burst_packed_ram_addr_269 = write_burst_packed_addr_259 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_270;
  assign write_burst_packed_ram_wdata_270 = _maxi_rdata_sb_0 >> 24;
  assign ram_w8_l16384_id1_3_1_wdata = ((write_burst_packed_fsm_13 == 1) && write_burst_block_ram_wvalid_257)? write_burst_packed_ram_wdata_270 : 'hx;
  assign ram_w8_l16384_id1_3_1_wenable = ((write_burst_packed_fsm_13 == 1) && write_burst_block_ram_wvalid_257)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_271;
  wire write_burst_block_ram_wquit_272;
  reg [32-1:0] write_burst_packed_fsm_14;
  localparam write_burst_packed_fsm_14_init = 0;
  reg [14-1:0] write_burst_packed_addr_273;
  reg [14-1:0] write_burst_packed_stride_274;
  reg [33-1:0] write_burst_packed_length_275;
  reg write_burst_packed_done_276;
  wire [12-1:0] write_burst_packed_ram_addr_277;
  assign write_burst_packed_ram_addr_277 = write_burst_packed_addr_273 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_278;
  assign write_burst_packed_ram_wdata_278 = _maxi_rdata_sb_0 >> 0;
  assign ram_w8_l16384_id2_0_1_addr = ((write_burst_packed_fsm_14 == 1) && write_burst_block_ram_wvalid_271)? write_burst_packed_ram_addr_277 : 'hx;
  assign ram_w8_l16384_id2_0_1_wdata = ((write_burst_packed_fsm_14 == 1) && write_burst_block_ram_wvalid_271)? write_burst_packed_ram_wdata_278 : 'hx;
  assign ram_w8_l16384_id2_0_1_wenable = ((write_burst_packed_fsm_14 == 1) && write_burst_block_ram_wvalid_271)? 1'd1 : 0;
  assign ram_w8_l16384_id2_0_1_enable = ((write_burst_packed_fsm_14 == 1) && write_burst_block_ram_wvalid_271)? 1'd1 : 0;
  wire [12-1:0] write_burst_packed_ram_addr_279;
  assign write_burst_packed_ram_addr_279 = write_burst_packed_addr_273 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_280;
  assign write_burst_packed_ram_wdata_280 = _maxi_rdata_sb_0 >> 8;
  assign ram_w8_l16384_id2_1_1_addr = ((write_burst_packed_fsm_14 == 1) && write_burst_block_ram_wvalid_271)? write_burst_packed_ram_addr_279 : 'hx;
  assign ram_w8_l16384_id2_1_1_wdata = ((write_burst_packed_fsm_14 == 1) && write_burst_block_ram_wvalid_271)? write_burst_packed_ram_wdata_280 : 'hx;
  assign ram_w8_l16384_id2_1_1_wenable = ((write_burst_packed_fsm_14 == 1) && write_burst_block_ram_wvalid_271)? 1'd1 : 0;
  assign ram_w8_l16384_id2_1_1_enable = ((write_burst_packed_fsm_14 == 1) && write_burst_block_ram_wvalid_271)? 1'd1 : 0;
  wire [12-1:0] write_burst_packed_ram_addr_281;
  assign write_burst_packed_ram_addr_281 = write_burst_packed_addr_273 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_282;
  assign write_burst_packed_ram_wdata_282 = _maxi_rdata_sb_0 >> 16;
  assign ram_w8_l16384_id2_2_1_addr = ((write_burst_packed_fsm_14 == 1) && write_burst_block_ram_wvalid_271)? write_burst_packed_ram_addr_281 : 'hx;
  assign ram_w8_l16384_id2_2_1_wdata = ((write_burst_packed_fsm_14 == 1) && write_burst_block_ram_wvalid_271)? write_burst_packed_ram_wdata_282 : 'hx;
  assign ram_w8_l16384_id2_2_1_wenable = ((write_burst_packed_fsm_14 == 1) && write_burst_block_ram_wvalid_271)? 1'd1 : 0;
  assign ram_w8_l16384_id2_2_1_enable = ((write_burst_packed_fsm_14 == 1) && write_burst_block_ram_wvalid_271)? 1'd1 : 0;
  wire [12-1:0] write_burst_packed_ram_addr_283;
  assign write_burst_packed_ram_addr_283 = write_burst_packed_addr_273 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_284;
  assign write_burst_packed_ram_wdata_284 = _maxi_rdata_sb_0 >> 24;
  assign ram_w8_l16384_id2_3_1_addr = ((write_burst_packed_fsm_14 == 1) && write_burst_block_ram_wvalid_271)? write_burst_packed_ram_addr_283 : 'hx;
  assign ram_w8_l16384_id2_3_1_wdata = ((write_burst_packed_fsm_14 == 1) && write_burst_block_ram_wvalid_271)? write_burst_packed_ram_wdata_284 : 'hx;
  assign ram_w8_l16384_id2_3_1_wenable = ((write_burst_packed_fsm_14 == 1) && write_burst_block_ram_wvalid_271)? 1'd1 : 0;
  assign ram_w8_l16384_id2_3_1_enable = ((write_burst_packed_fsm_14 == 1) && write_burst_block_ram_wvalid_271)? 1'd1 : 0;
  reg [32-1:0] write_burst_block_fsm_15;
  localparam write_burst_block_fsm_15_init = 0;
  reg [33-1:0] write_burst_block_length_285;
  reg [32-1:0] write_burst_block_blocksize_286;
  reg write_burst_block_done_287;
  reg [32-1:0] write_burst_block_count_288;
  assign write_burst_block_ram_wvalid_243 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_15 == 1);
  assign write_burst_block_ram_wquit_244 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_285 <= 1);
  assign write_burst_block_ram_wvalid_257 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_15 == 2);
  assign write_burst_block_ram_wquit_258 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_285 <= 1);
  assign write_burst_block_ram_wvalid_271 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_15 == 3);
  assign write_burst_block_ram_wquit_272 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_285 <= 1);
  wire [14-1:0] _dma_write_block_high_local_size_289;
  assign _dma_write_block_high_local_size_289 = cparam_conv2d_24_act_read_size >> 2;
  wire [2-1:0] _dma_write_block_low_local_size_290;
  assign _dma_write_block_low_local_size_290 = cparam_conv2d_24_act_read_size & { 2{ 1'd1 } };
  wire [14-1:0] _dma_write_block_local_size_291;
  assign _dma_write_block_local_size_291 = (_dma_write_block_low_local_size_290 > 0)? _dma_write_block_high_local_size_289 + 1 : _dma_write_block_high_local_size_289;
  wire [10-1:0] _dma_read_block_high_local_blocksize_292;
  assign _dma_read_block_high_local_blocksize_292 = cparam_conv2d_24_act_read_block >> 2;
  wire [3-1:0] _dma_read_block_low_local_blocksize_293;
  assign _dma_read_block_low_local_blocksize_293 = cparam_conv2d_24_act_read_block & { 2{ 1'd1 } };
  wire [10-1:0] _dma_read_block_local_blocksize_294;
  assign _dma_read_block_local_blocksize_294 = (_dma_read_block_low_local_blocksize_293 > 0)? _dma_read_block_high_local_blocksize_292 + 1 : _dma_read_block_high_local_blocksize_292;
  wire [32-1:0] mask_addr_shifted_295;
  assign mask_addr_shifted_295 = conv2d_24_mux_act_gaddr_1 + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_296;
  assign mask_addr_masked_296 = mask_addr_shifted_295 << 2;
  wire write_burst_block_ram_wvalid_297;
  wire write_burst_block_ram_wquit_298;
  reg [32-1:0] write_burst_packed_fsm_16;
  localparam write_burst_packed_fsm_16_init = 0;
  reg [14-1:0] write_burst_packed_addr_299;
  reg [14-1:0] write_burst_packed_stride_300;
  reg [33-1:0] write_burst_packed_length_301;
  reg write_burst_packed_done_302;
  wire [12-1:0] write_burst_packed_ram_addr_303;
  assign write_burst_packed_ram_addr_303 = write_burst_packed_addr_299 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_304;
  assign write_burst_packed_ram_wdata_304 = _maxi_rdata_sb_0 >> 0;
  assign ram_w8_l16384_id3_0_1_addr = ((write_burst_packed_fsm_16 == 1) && write_burst_block_ram_wvalid_297)? write_burst_packed_ram_addr_303 : 'hx;
  assign ram_w8_l16384_id3_0_1_wdata = ((write_burst_packed_fsm_16 == 1) && write_burst_block_ram_wvalid_297)? write_burst_packed_ram_wdata_304 : 'hx;
  assign ram_w8_l16384_id3_0_1_wenable = ((write_burst_packed_fsm_16 == 1) && write_burst_block_ram_wvalid_297)? 1'd1 : 0;
  assign ram_w8_l16384_id3_0_1_enable = ((write_burst_packed_fsm_16 == 1) && write_burst_block_ram_wvalid_297)? 1'd1 : 0;
  wire [12-1:0] write_burst_packed_ram_addr_305;
  assign write_burst_packed_ram_addr_305 = write_burst_packed_addr_299 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_306;
  assign write_burst_packed_ram_wdata_306 = _maxi_rdata_sb_0 >> 8;
  assign ram_w8_l16384_id3_1_1_addr = ((write_burst_packed_fsm_16 == 1) && write_burst_block_ram_wvalid_297)? write_burst_packed_ram_addr_305 : 'hx;
  assign ram_w8_l16384_id3_1_1_wdata = ((write_burst_packed_fsm_16 == 1) && write_burst_block_ram_wvalid_297)? write_burst_packed_ram_wdata_306 : 'hx;
  assign ram_w8_l16384_id3_1_1_wenable = ((write_burst_packed_fsm_16 == 1) && write_burst_block_ram_wvalid_297)? 1'd1 : 0;
  assign ram_w8_l16384_id3_1_1_enable = ((write_burst_packed_fsm_16 == 1) && write_burst_block_ram_wvalid_297)? 1'd1 : 0;
  wire [12-1:0] write_burst_packed_ram_addr_307;
  assign write_burst_packed_ram_addr_307 = write_burst_packed_addr_299 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_308;
  assign write_burst_packed_ram_wdata_308 = _maxi_rdata_sb_0 >> 16;
  assign ram_w8_l16384_id3_2_1_addr = ((write_burst_packed_fsm_16 == 1) && write_burst_block_ram_wvalid_297)? write_burst_packed_ram_addr_307 : 'hx;
  assign ram_w8_l16384_id3_2_1_wdata = ((write_burst_packed_fsm_16 == 1) && write_burst_block_ram_wvalid_297)? write_burst_packed_ram_wdata_308 : 'hx;
  assign ram_w8_l16384_id3_2_1_wenable = ((write_burst_packed_fsm_16 == 1) && write_burst_block_ram_wvalid_297)? 1'd1 : 0;
  assign ram_w8_l16384_id3_2_1_enable = ((write_burst_packed_fsm_16 == 1) && write_burst_block_ram_wvalid_297)? 1'd1 : 0;
  wire [12-1:0] write_burst_packed_ram_addr_309;
  assign write_burst_packed_ram_addr_309 = write_burst_packed_addr_299 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_310;
  assign write_burst_packed_ram_wdata_310 = _maxi_rdata_sb_0 >> 24;
  assign ram_w8_l16384_id3_3_1_addr = ((write_burst_packed_fsm_16 == 1) && write_burst_block_ram_wvalid_297)? write_burst_packed_ram_addr_309 : 'hx;
  assign ram_w8_l16384_id3_3_1_wdata = ((write_burst_packed_fsm_16 == 1) && write_burst_block_ram_wvalid_297)? write_burst_packed_ram_wdata_310 : 'hx;
  assign ram_w8_l16384_id3_3_1_wenable = ((write_burst_packed_fsm_16 == 1) && write_burst_block_ram_wvalid_297)? 1'd1 : 0;
  assign ram_w8_l16384_id3_3_1_enable = ((write_burst_packed_fsm_16 == 1) && write_burst_block_ram_wvalid_297)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_311;
  wire write_burst_block_ram_wquit_312;
  reg [32-1:0] write_burst_packed_fsm_17;
  localparam write_burst_packed_fsm_17_init = 0;
  reg [14-1:0] write_burst_packed_addr_313;
  reg [14-1:0] write_burst_packed_stride_314;
  reg [33-1:0] write_burst_packed_length_315;
  reg write_burst_packed_done_316;
  wire [12-1:0] write_burst_packed_ram_addr_317;
  assign write_burst_packed_ram_addr_317 = write_burst_packed_addr_313 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_318;
  assign write_burst_packed_ram_wdata_318 = _maxi_rdata_sb_0 >> 0;
  assign ram_w8_l16384_id4_0_1_addr = ((write_burst_packed_fsm_17 == 1) && write_burst_block_ram_wvalid_311)? write_burst_packed_ram_addr_317 : 'hx;
  assign ram_w8_l16384_id4_0_1_wdata = ((write_burst_packed_fsm_17 == 1) && write_burst_block_ram_wvalid_311)? write_burst_packed_ram_wdata_318 : 'hx;
  assign ram_w8_l16384_id4_0_1_wenable = ((write_burst_packed_fsm_17 == 1) && write_burst_block_ram_wvalid_311)? 1'd1 : 0;
  assign ram_w8_l16384_id4_0_1_enable = ((write_burst_packed_fsm_17 == 1) && write_burst_block_ram_wvalid_311)? 1'd1 : 0;
  wire [12-1:0] write_burst_packed_ram_addr_319;
  assign write_burst_packed_ram_addr_319 = write_burst_packed_addr_313 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_320;
  assign write_burst_packed_ram_wdata_320 = _maxi_rdata_sb_0 >> 8;
  assign ram_w8_l16384_id4_1_1_addr = ((write_burst_packed_fsm_17 == 1) && write_burst_block_ram_wvalid_311)? write_burst_packed_ram_addr_319 : 'hx;
  assign ram_w8_l16384_id4_1_1_wdata = ((write_burst_packed_fsm_17 == 1) && write_burst_block_ram_wvalid_311)? write_burst_packed_ram_wdata_320 : 'hx;
  assign ram_w8_l16384_id4_1_1_wenable = ((write_burst_packed_fsm_17 == 1) && write_burst_block_ram_wvalid_311)? 1'd1 : 0;
  assign ram_w8_l16384_id4_1_1_enable = ((write_burst_packed_fsm_17 == 1) && write_burst_block_ram_wvalid_311)? 1'd1 : 0;
  wire [12-1:0] write_burst_packed_ram_addr_321;
  assign write_burst_packed_ram_addr_321 = write_burst_packed_addr_313 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_322;
  assign write_burst_packed_ram_wdata_322 = _maxi_rdata_sb_0 >> 16;
  assign ram_w8_l16384_id4_2_1_addr = ((write_burst_packed_fsm_17 == 1) && write_burst_block_ram_wvalid_311)? write_burst_packed_ram_addr_321 : 'hx;
  assign ram_w8_l16384_id4_2_1_wdata = ((write_burst_packed_fsm_17 == 1) && write_burst_block_ram_wvalid_311)? write_burst_packed_ram_wdata_322 : 'hx;
  assign ram_w8_l16384_id4_2_1_wenable = ((write_burst_packed_fsm_17 == 1) && write_burst_block_ram_wvalid_311)? 1'd1 : 0;
  assign ram_w8_l16384_id4_2_1_enable = ((write_burst_packed_fsm_17 == 1) && write_burst_block_ram_wvalid_311)? 1'd1 : 0;
  wire [12-1:0] write_burst_packed_ram_addr_323;
  assign write_burst_packed_ram_addr_323 = write_burst_packed_addr_313 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_324;
  assign write_burst_packed_ram_wdata_324 = _maxi_rdata_sb_0 >> 24;
  assign ram_w8_l16384_id4_3_1_addr = ((write_burst_packed_fsm_17 == 1) && write_burst_block_ram_wvalid_311)? write_burst_packed_ram_addr_323 : 'hx;
  assign ram_w8_l16384_id4_3_1_wdata = ((write_burst_packed_fsm_17 == 1) && write_burst_block_ram_wvalid_311)? write_burst_packed_ram_wdata_324 : 'hx;
  assign ram_w8_l16384_id4_3_1_wenable = ((write_burst_packed_fsm_17 == 1) && write_burst_block_ram_wvalid_311)? 1'd1 : 0;
  assign ram_w8_l16384_id4_3_1_enable = ((write_burst_packed_fsm_17 == 1) && write_burst_block_ram_wvalid_311)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_325;
  wire write_burst_block_ram_wquit_326;
  reg [32-1:0] write_burst_packed_fsm_18;
  localparam write_burst_packed_fsm_18_init = 0;
  reg [14-1:0] write_burst_packed_addr_327;
  reg [14-1:0] write_burst_packed_stride_328;
  reg [33-1:0] write_burst_packed_length_329;
  reg write_burst_packed_done_330;
  wire [12-1:0] write_burst_packed_ram_addr_331;
  assign write_burst_packed_ram_addr_331 = write_burst_packed_addr_327 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_332;
  assign write_burst_packed_ram_wdata_332 = _maxi_rdata_sb_0 >> 0;
  assign ram_w8_l16384_id5_0_1_addr = ((write_burst_packed_fsm_18 == 1) && write_burst_block_ram_wvalid_325)? write_burst_packed_ram_addr_331 : 'hx;
  assign ram_w8_l16384_id5_0_1_wdata = ((write_burst_packed_fsm_18 == 1) && write_burst_block_ram_wvalid_325)? write_burst_packed_ram_wdata_332 : 'hx;
  assign ram_w8_l16384_id5_0_1_wenable = ((write_burst_packed_fsm_18 == 1) && write_burst_block_ram_wvalid_325)? 1'd1 : 0;
  assign ram_w8_l16384_id5_0_1_enable = ((write_burst_packed_fsm_18 == 1) && write_burst_block_ram_wvalid_325)? 1'd1 : 0;
  wire [12-1:0] write_burst_packed_ram_addr_333;
  assign write_burst_packed_ram_addr_333 = write_burst_packed_addr_327 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_334;
  assign write_burst_packed_ram_wdata_334 = _maxi_rdata_sb_0 >> 8;
  assign ram_w8_l16384_id5_1_1_addr = ((write_burst_packed_fsm_18 == 1) && write_burst_block_ram_wvalid_325)? write_burst_packed_ram_addr_333 : 'hx;
  assign ram_w8_l16384_id5_1_1_wdata = ((write_burst_packed_fsm_18 == 1) && write_burst_block_ram_wvalid_325)? write_burst_packed_ram_wdata_334 : 'hx;
  assign ram_w8_l16384_id5_1_1_wenable = ((write_burst_packed_fsm_18 == 1) && write_burst_block_ram_wvalid_325)? 1'd1 : 0;
  assign ram_w8_l16384_id5_1_1_enable = ((write_burst_packed_fsm_18 == 1) && write_burst_block_ram_wvalid_325)? 1'd1 : 0;
  wire [12-1:0] write_burst_packed_ram_addr_335;
  assign write_burst_packed_ram_addr_335 = write_burst_packed_addr_327 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_336;
  assign write_burst_packed_ram_wdata_336 = _maxi_rdata_sb_0 >> 16;
  assign ram_w8_l16384_id5_2_1_addr = ((write_burst_packed_fsm_18 == 1) && write_burst_block_ram_wvalid_325)? write_burst_packed_ram_addr_335 : 'hx;
  assign ram_w8_l16384_id5_2_1_wdata = ((write_burst_packed_fsm_18 == 1) && write_burst_block_ram_wvalid_325)? write_burst_packed_ram_wdata_336 : 'hx;
  assign ram_w8_l16384_id5_2_1_wenable = ((write_burst_packed_fsm_18 == 1) && write_burst_block_ram_wvalid_325)? 1'd1 : 0;
  assign ram_w8_l16384_id5_2_1_enable = ((write_burst_packed_fsm_18 == 1) && write_burst_block_ram_wvalid_325)? 1'd1 : 0;
  wire [12-1:0] write_burst_packed_ram_addr_337;
  assign write_burst_packed_ram_addr_337 = write_burst_packed_addr_327 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_338;
  assign write_burst_packed_ram_wdata_338 = _maxi_rdata_sb_0 >> 24;
  assign ram_w8_l16384_id5_3_1_addr = ((write_burst_packed_fsm_18 == 1) && write_burst_block_ram_wvalid_325)? write_burst_packed_ram_addr_337 : 'hx;
  assign ram_w8_l16384_id5_3_1_wdata = ((write_burst_packed_fsm_18 == 1) && write_burst_block_ram_wvalid_325)? write_burst_packed_ram_wdata_338 : 'hx;
  assign ram_w8_l16384_id5_3_1_wenable = ((write_burst_packed_fsm_18 == 1) && write_burst_block_ram_wvalid_325)? 1'd1 : 0;
  assign ram_w8_l16384_id5_3_1_enable = ((write_burst_packed_fsm_18 == 1) && write_burst_block_ram_wvalid_325)? 1'd1 : 0;
  reg [32-1:0] write_burst_block_fsm_19;
  localparam write_burst_block_fsm_19_init = 0;
  reg [33-1:0] write_burst_block_length_339;
  reg [32-1:0] write_burst_block_blocksize_340;
  reg write_burst_block_done_341;
  reg [32-1:0] write_burst_block_count_342;
  assign write_burst_block_ram_wvalid_297 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_19 == 1);
  assign write_burst_block_ram_wquit_298 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_339 <= 1);
  assign write_burst_block_ram_wvalid_311 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_19 == 2);
  assign write_burst_block_ram_wquit_312 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_339 <= 1);
  assign write_burst_block_ram_wvalid_325 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_19 == 3);
  assign write_burst_block_ram_wquit_326 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_339 <= 1);
  wire [14-1:0] _dma_write_block_high_local_size_343;
  assign _dma_write_block_high_local_size_343 = cparam_conv2d_24_act_read_size >> 2;
  wire [2-1:0] _dma_write_block_low_local_size_344;
  assign _dma_write_block_low_local_size_344 = cparam_conv2d_24_act_read_size & { 2{ 1'd1 } };
  wire [14-1:0] _dma_write_block_local_size_345;
  assign _dma_write_block_local_size_345 = (_dma_write_block_low_local_size_344 > 0)? _dma_write_block_high_local_size_343 + 1 : _dma_write_block_high_local_size_343;
  wire [10-1:0] _dma_read_block_high_local_blocksize_346;
  assign _dma_read_block_high_local_blocksize_346 = cparam_conv2d_24_act_read_block >> 2;
  wire [3-1:0] _dma_read_block_low_local_blocksize_347;
  assign _dma_read_block_low_local_blocksize_347 = cparam_conv2d_24_act_read_block & { 2{ 1'd1 } };
  wire [10-1:0] _dma_read_block_local_blocksize_348;
  assign _dma_read_block_local_blocksize_348 = (_dma_read_block_low_local_blocksize_347 > 0)? _dma_read_block_high_local_blocksize_346 + 1 : _dma_read_block_high_local_blocksize_346;
  wire [32-1:0] mask_addr_shifted_349;
  assign mask_addr_shifted_349 = conv2d_24_mux_act_gaddr_2 + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_350;
  assign mask_addr_masked_350 = mask_addr_shifted_349 << 2;
  wire write_burst_block_ram_wvalid_351;
  wire write_burst_block_ram_wquit_352;
  reg [32-1:0] write_burst_packed_fsm_20;
  localparam write_burst_packed_fsm_20_init = 0;
  reg [14-1:0] write_burst_packed_addr_353;
  reg [14-1:0] write_burst_packed_stride_354;
  reg [33-1:0] write_burst_packed_length_355;
  reg write_burst_packed_done_356;
  wire [12-1:0] write_burst_packed_ram_addr_357;
  assign write_burst_packed_ram_addr_357 = write_burst_packed_addr_353 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_358;
  assign write_burst_packed_ram_wdata_358 = _maxi_rdata_sb_0 >> 0;
  assign ram_w8_l16384_id6_0_1_addr = ((write_burst_packed_fsm_20 == 1) && write_burst_block_ram_wvalid_351)? write_burst_packed_ram_addr_357 : 'hx;
  assign ram_w8_l16384_id6_0_1_wdata = ((write_burst_packed_fsm_20 == 1) && write_burst_block_ram_wvalid_351)? write_burst_packed_ram_wdata_358 : 'hx;
  assign ram_w8_l16384_id6_0_1_wenable = ((write_burst_packed_fsm_20 == 1) && write_burst_block_ram_wvalid_351)? 1'd1 : 0;
  assign ram_w8_l16384_id6_0_1_enable = ((write_burst_packed_fsm_20 == 1) && write_burst_block_ram_wvalid_351)? 1'd1 : 0;
  wire [12-1:0] write_burst_packed_ram_addr_359;
  assign write_burst_packed_ram_addr_359 = write_burst_packed_addr_353 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_360;
  assign write_burst_packed_ram_wdata_360 = _maxi_rdata_sb_0 >> 8;
  assign ram_w8_l16384_id6_1_1_addr = ((write_burst_packed_fsm_20 == 1) && write_burst_block_ram_wvalid_351)? write_burst_packed_ram_addr_359 : 'hx;
  assign ram_w8_l16384_id6_1_1_wdata = ((write_burst_packed_fsm_20 == 1) && write_burst_block_ram_wvalid_351)? write_burst_packed_ram_wdata_360 : 'hx;
  assign ram_w8_l16384_id6_1_1_wenable = ((write_burst_packed_fsm_20 == 1) && write_burst_block_ram_wvalid_351)? 1'd1 : 0;
  assign ram_w8_l16384_id6_1_1_enable = ((write_burst_packed_fsm_20 == 1) && write_burst_block_ram_wvalid_351)? 1'd1 : 0;
  wire [12-1:0] write_burst_packed_ram_addr_361;
  assign write_burst_packed_ram_addr_361 = write_burst_packed_addr_353 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_362;
  assign write_burst_packed_ram_wdata_362 = _maxi_rdata_sb_0 >> 16;
  assign ram_w8_l16384_id6_2_1_addr = ((write_burst_packed_fsm_20 == 1) && write_burst_block_ram_wvalid_351)? write_burst_packed_ram_addr_361 : 'hx;
  assign ram_w8_l16384_id6_2_1_wdata = ((write_burst_packed_fsm_20 == 1) && write_burst_block_ram_wvalid_351)? write_burst_packed_ram_wdata_362 : 'hx;
  assign ram_w8_l16384_id6_2_1_wenable = ((write_burst_packed_fsm_20 == 1) && write_burst_block_ram_wvalid_351)? 1'd1 : 0;
  assign ram_w8_l16384_id6_2_1_enable = ((write_burst_packed_fsm_20 == 1) && write_burst_block_ram_wvalid_351)? 1'd1 : 0;
  wire [12-1:0] write_burst_packed_ram_addr_363;
  assign write_burst_packed_ram_addr_363 = write_burst_packed_addr_353 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_364;
  assign write_burst_packed_ram_wdata_364 = _maxi_rdata_sb_0 >> 24;
  assign ram_w8_l16384_id6_3_1_addr = ((write_burst_packed_fsm_20 == 1) && write_burst_block_ram_wvalid_351)? write_burst_packed_ram_addr_363 : 'hx;
  assign ram_w8_l16384_id6_3_1_wdata = ((write_burst_packed_fsm_20 == 1) && write_burst_block_ram_wvalid_351)? write_burst_packed_ram_wdata_364 : 'hx;
  assign ram_w8_l16384_id6_3_1_wenable = ((write_burst_packed_fsm_20 == 1) && write_burst_block_ram_wvalid_351)? 1'd1 : 0;
  assign ram_w8_l16384_id6_3_1_enable = ((write_burst_packed_fsm_20 == 1) && write_burst_block_ram_wvalid_351)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_365;
  wire write_burst_block_ram_wquit_366;
  reg [32-1:0] write_burst_packed_fsm_21;
  localparam write_burst_packed_fsm_21_init = 0;
  reg [14-1:0] write_burst_packed_addr_367;
  reg [14-1:0] write_burst_packed_stride_368;
  reg [33-1:0] write_burst_packed_length_369;
  reg write_burst_packed_done_370;
  wire [12-1:0] write_burst_packed_ram_addr_371;
  assign write_burst_packed_ram_addr_371 = write_burst_packed_addr_367 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_372;
  assign write_burst_packed_ram_wdata_372 = _maxi_rdata_sb_0 >> 0;
  assign ram_w8_l16384_id7_0_1_addr = ((write_burst_packed_fsm_21 == 1) && write_burst_block_ram_wvalid_365)? write_burst_packed_ram_addr_371 : 'hx;
  assign ram_w8_l16384_id7_0_1_wdata = ((write_burst_packed_fsm_21 == 1) && write_burst_block_ram_wvalid_365)? write_burst_packed_ram_wdata_372 : 'hx;
  assign ram_w8_l16384_id7_0_1_wenable = ((write_burst_packed_fsm_21 == 1) && write_burst_block_ram_wvalid_365)? 1'd1 : 0;
  assign ram_w8_l16384_id7_0_1_enable = ((write_burst_packed_fsm_21 == 1) && write_burst_block_ram_wvalid_365)? 1'd1 : 0;
  wire [12-1:0] write_burst_packed_ram_addr_373;
  assign write_burst_packed_ram_addr_373 = write_burst_packed_addr_367 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_374;
  assign write_burst_packed_ram_wdata_374 = _maxi_rdata_sb_0 >> 8;
  assign ram_w8_l16384_id7_1_1_addr = ((write_burst_packed_fsm_21 == 1) && write_burst_block_ram_wvalid_365)? write_burst_packed_ram_addr_373 : 'hx;
  assign ram_w8_l16384_id7_1_1_wdata = ((write_burst_packed_fsm_21 == 1) && write_burst_block_ram_wvalid_365)? write_burst_packed_ram_wdata_374 : 'hx;
  assign ram_w8_l16384_id7_1_1_wenable = ((write_burst_packed_fsm_21 == 1) && write_burst_block_ram_wvalid_365)? 1'd1 : 0;
  assign ram_w8_l16384_id7_1_1_enable = ((write_burst_packed_fsm_21 == 1) && write_burst_block_ram_wvalid_365)? 1'd1 : 0;
  wire [12-1:0] write_burst_packed_ram_addr_375;
  assign write_burst_packed_ram_addr_375 = write_burst_packed_addr_367 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_376;
  assign write_burst_packed_ram_wdata_376 = _maxi_rdata_sb_0 >> 16;
  assign ram_w8_l16384_id7_2_1_addr = ((write_burst_packed_fsm_21 == 1) && write_burst_block_ram_wvalid_365)? write_burst_packed_ram_addr_375 : 'hx;
  assign ram_w8_l16384_id7_2_1_wdata = ((write_burst_packed_fsm_21 == 1) && write_burst_block_ram_wvalid_365)? write_burst_packed_ram_wdata_376 : 'hx;
  assign ram_w8_l16384_id7_2_1_wenable = ((write_burst_packed_fsm_21 == 1) && write_burst_block_ram_wvalid_365)? 1'd1 : 0;
  assign ram_w8_l16384_id7_2_1_enable = ((write_burst_packed_fsm_21 == 1) && write_burst_block_ram_wvalid_365)? 1'd1 : 0;
  wire [12-1:0] write_burst_packed_ram_addr_377;
  assign write_burst_packed_ram_addr_377 = write_burst_packed_addr_367 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_378;
  assign write_burst_packed_ram_wdata_378 = _maxi_rdata_sb_0 >> 24;
  assign ram_w8_l16384_id7_3_1_addr = ((write_burst_packed_fsm_21 == 1) && write_burst_block_ram_wvalid_365)? write_burst_packed_ram_addr_377 : 'hx;
  assign ram_w8_l16384_id7_3_1_wdata = ((write_burst_packed_fsm_21 == 1) && write_burst_block_ram_wvalid_365)? write_burst_packed_ram_wdata_378 : 'hx;
  assign ram_w8_l16384_id7_3_1_wenable = ((write_burst_packed_fsm_21 == 1) && write_burst_block_ram_wvalid_365)? 1'd1 : 0;
  assign ram_w8_l16384_id7_3_1_enable = ((write_burst_packed_fsm_21 == 1) && write_burst_block_ram_wvalid_365)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_379;
  wire write_burst_block_ram_wquit_380;
  reg [32-1:0] write_burst_packed_fsm_22;
  localparam write_burst_packed_fsm_22_init = 0;
  reg [14-1:0] write_burst_packed_addr_381;
  reg [14-1:0] write_burst_packed_stride_382;
  reg [33-1:0] write_burst_packed_length_383;
  reg write_burst_packed_done_384;
  wire [12-1:0] write_burst_packed_ram_addr_385;
  assign write_burst_packed_ram_addr_385 = write_burst_packed_addr_381 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_386;
  assign write_burst_packed_ram_wdata_386 = _maxi_rdata_sb_0 >> 0;
  assign ram_w8_l16384_id8_0_1_addr = ((write_burst_packed_fsm_22 == 1) && write_burst_block_ram_wvalid_379)? write_burst_packed_ram_addr_385 : 'hx;
  assign ram_w8_l16384_id8_0_1_wdata = ((write_burst_packed_fsm_22 == 1) && write_burst_block_ram_wvalid_379)? write_burst_packed_ram_wdata_386 : 'hx;
  assign ram_w8_l16384_id8_0_1_wenable = ((write_burst_packed_fsm_22 == 1) && write_burst_block_ram_wvalid_379)? 1'd1 : 0;
  assign ram_w8_l16384_id8_0_1_enable = ((write_burst_packed_fsm_22 == 1) && write_burst_block_ram_wvalid_379)? 1'd1 : 0;
  wire [12-1:0] write_burst_packed_ram_addr_387;
  assign write_burst_packed_ram_addr_387 = write_burst_packed_addr_381 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_388;
  assign write_burst_packed_ram_wdata_388 = _maxi_rdata_sb_0 >> 8;
  assign ram_w8_l16384_id8_1_1_addr = ((write_burst_packed_fsm_22 == 1) && write_burst_block_ram_wvalid_379)? write_burst_packed_ram_addr_387 : 'hx;
  assign ram_w8_l16384_id8_1_1_wdata = ((write_burst_packed_fsm_22 == 1) && write_burst_block_ram_wvalid_379)? write_burst_packed_ram_wdata_388 : 'hx;
  assign ram_w8_l16384_id8_1_1_wenable = ((write_burst_packed_fsm_22 == 1) && write_burst_block_ram_wvalid_379)? 1'd1 : 0;
  assign ram_w8_l16384_id8_1_1_enable = ((write_burst_packed_fsm_22 == 1) && write_burst_block_ram_wvalid_379)? 1'd1 : 0;
  wire [12-1:0] write_burst_packed_ram_addr_389;
  assign write_burst_packed_ram_addr_389 = write_burst_packed_addr_381 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_390;
  assign write_burst_packed_ram_wdata_390 = _maxi_rdata_sb_0 >> 16;
  assign ram_w8_l16384_id8_2_1_addr = ((write_burst_packed_fsm_22 == 1) && write_burst_block_ram_wvalid_379)? write_burst_packed_ram_addr_389 : 'hx;
  assign ram_w8_l16384_id8_2_1_wdata = ((write_burst_packed_fsm_22 == 1) && write_burst_block_ram_wvalid_379)? write_burst_packed_ram_wdata_390 : 'hx;
  assign ram_w8_l16384_id8_2_1_wenable = ((write_burst_packed_fsm_22 == 1) && write_burst_block_ram_wvalid_379)? 1'd1 : 0;
  assign ram_w8_l16384_id8_2_1_enable = ((write_burst_packed_fsm_22 == 1) && write_burst_block_ram_wvalid_379)? 1'd1 : 0;
  wire [12-1:0] write_burst_packed_ram_addr_391;
  assign write_burst_packed_ram_addr_391 = write_burst_packed_addr_381 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_392;
  assign write_burst_packed_ram_wdata_392 = _maxi_rdata_sb_0 >> 24;
  assign ram_w8_l16384_id8_3_1_addr = ((write_burst_packed_fsm_22 == 1) && write_burst_block_ram_wvalid_379)? write_burst_packed_ram_addr_391 : 'hx;
  assign ram_w8_l16384_id8_3_1_wdata = ((write_burst_packed_fsm_22 == 1) && write_burst_block_ram_wvalid_379)? write_burst_packed_ram_wdata_392 : 'hx;
  assign ram_w8_l16384_id8_3_1_wenable = ((write_burst_packed_fsm_22 == 1) && write_burst_block_ram_wvalid_379)? 1'd1 : 0;
  assign ram_w8_l16384_id8_3_1_enable = ((write_burst_packed_fsm_22 == 1) && write_burst_block_ram_wvalid_379)? 1'd1 : 0;
  reg [32-1:0] write_burst_block_fsm_23;
  localparam write_burst_block_fsm_23_init = 0;
  reg [33-1:0] write_burst_block_length_393;
  reg [32-1:0] write_burst_block_blocksize_394;
  reg write_burst_block_done_395;
  reg [32-1:0] write_burst_block_count_396;
  assign write_burst_block_ram_wvalid_351 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_23 == 1);
  assign write_burst_block_ram_wquit_352 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_393 <= 1);
  assign write_burst_block_ram_wvalid_365 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_23 == 2);
  assign write_burst_block_ram_wquit_366 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_393 <= 1);
  assign write_burst_block_ram_wvalid_379 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_23 == 3);
  assign write_burst_block_ram_wquit_380 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_393 <= 1);
  reg [32-1:0] conv2d_24_comp_fsm;
  localparam conv2d_24_comp_fsm_init = 0;
  reg [32-1:0] conv2d_24_filter_page_comp_offset_buf;
  reg [32-1:0] conv2d_24_act_page_comp_offset_buf_0;
  reg [32-1:0] conv2d_24_act_page_comp_offset_buf_1;
  reg [32-1:0] conv2d_24_act_page_comp_offset_buf_2;
  reg [32-1:0] conv2d_24_out_page_comp_offset_buf;
  reg [32-1:0] conv2d_24_row_count_buf;
  reg [2-1:0] conv2d_24_row_select_buf;
  reg [32-1:0] conv2d_24_och_count_buf;
  wire conv2d_24_stream_pad_mask_0_0;
  assign conv2d_24_stream_pad_mask_0_0 = (conv2d_24_col_count + 0 < cparam_conv2d_24_pad_col_left) || (conv2d_24_col_count + 0 >= cparam_conv2d_24_act_num_col + cparam_conv2d_24_pad_col_left) || (conv2d_24_row_count_buf + 0 < cparam_conv2d_24_pad_row_top) || (conv2d_24_row_count_buf + 0 >= cparam_conv2d_24_act_num_row + cparam_conv2d_24_pad_row_top);
  wire conv2d_24_stream_pad_mask_0_1;
  assign conv2d_24_stream_pad_mask_0_1 = (conv2d_24_col_count + 1 < cparam_conv2d_24_pad_col_left) || (conv2d_24_col_count + 1 >= cparam_conv2d_24_act_num_col + cparam_conv2d_24_pad_col_left) || (conv2d_24_row_count_buf + 0 < cparam_conv2d_24_pad_row_top) || (conv2d_24_row_count_buf + 0 >= cparam_conv2d_24_act_num_row + cparam_conv2d_24_pad_row_top);
  wire conv2d_24_stream_pad_mask_0_2;
  assign conv2d_24_stream_pad_mask_0_2 = (conv2d_24_col_count + 2 < cparam_conv2d_24_pad_col_left) || (conv2d_24_col_count + 2 >= cparam_conv2d_24_act_num_col + cparam_conv2d_24_pad_col_left) || (conv2d_24_row_count_buf + 0 < cparam_conv2d_24_pad_row_top) || (conv2d_24_row_count_buf + 0 >= cparam_conv2d_24_act_num_row + cparam_conv2d_24_pad_row_top);
  wire conv2d_24_stream_pad_mask_1_0;
  assign conv2d_24_stream_pad_mask_1_0 = (conv2d_24_col_count + 0 < cparam_conv2d_24_pad_col_left) || (conv2d_24_col_count + 0 >= cparam_conv2d_24_act_num_col + cparam_conv2d_24_pad_col_left) || (conv2d_24_row_count_buf + 1 < cparam_conv2d_24_pad_row_top) || (conv2d_24_row_count_buf + 1 >= cparam_conv2d_24_act_num_row + cparam_conv2d_24_pad_row_top);
  wire conv2d_24_stream_pad_mask_1_1;
  assign conv2d_24_stream_pad_mask_1_1 = (conv2d_24_col_count + 1 < cparam_conv2d_24_pad_col_left) || (conv2d_24_col_count + 1 >= cparam_conv2d_24_act_num_col + cparam_conv2d_24_pad_col_left) || (conv2d_24_row_count_buf + 1 < cparam_conv2d_24_pad_row_top) || (conv2d_24_row_count_buf + 1 >= cparam_conv2d_24_act_num_row + cparam_conv2d_24_pad_row_top);
  wire conv2d_24_stream_pad_mask_1_2;
  assign conv2d_24_stream_pad_mask_1_2 = (conv2d_24_col_count + 2 < cparam_conv2d_24_pad_col_left) || (conv2d_24_col_count + 2 >= cparam_conv2d_24_act_num_col + cparam_conv2d_24_pad_col_left) || (conv2d_24_row_count_buf + 1 < cparam_conv2d_24_pad_row_top) || (conv2d_24_row_count_buf + 1 >= cparam_conv2d_24_act_num_row + cparam_conv2d_24_pad_row_top);
  wire conv2d_24_stream_pad_mask_2_0;
  assign conv2d_24_stream_pad_mask_2_0 = (conv2d_24_col_count + 0 < cparam_conv2d_24_pad_col_left) || (conv2d_24_col_count + 0 >= cparam_conv2d_24_act_num_col + cparam_conv2d_24_pad_col_left) || (conv2d_24_row_count_buf + 2 < cparam_conv2d_24_pad_row_top) || (conv2d_24_row_count_buf + 2 >= cparam_conv2d_24_act_num_row + cparam_conv2d_24_pad_row_top);
  wire conv2d_24_stream_pad_mask_2_1;
  assign conv2d_24_stream_pad_mask_2_1 = (conv2d_24_col_count + 1 < cparam_conv2d_24_pad_col_left) || (conv2d_24_col_count + 1 >= cparam_conv2d_24_act_num_col + cparam_conv2d_24_pad_col_left) || (conv2d_24_row_count_buf + 2 < cparam_conv2d_24_pad_row_top) || (conv2d_24_row_count_buf + 2 >= cparam_conv2d_24_act_num_row + cparam_conv2d_24_pad_row_top);
  wire conv2d_24_stream_pad_mask_2_2;
  assign conv2d_24_stream_pad_mask_2_2 = (conv2d_24_col_count + 2 < cparam_conv2d_24_pad_col_left) || (conv2d_24_col_count + 2 >= cparam_conv2d_24_act_num_col + cparam_conv2d_24_pad_col_left) || (conv2d_24_row_count_buf + 2 < cparam_conv2d_24_pad_row_top) || (conv2d_24_row_count_buf + 2 >= cparam_conv2d_24_act_num_row + cparam_conv2d_24_pad_row_top);
  reg [9-1:0] conv2d_24_stream_pad_masks;
  wire [10-1:0] stream_conv2d_24_parameter_0_data;
  wire [2-1:0] stream_conv2d_24_parameter_1_data;
  wire [2-1:0] stream_conv2d_24_parameter_2_data;
  wire [9-1:0] stream_conv2d_24_parameter_3_data;
  wire [1-1:0] stream_conv2d_24_parameter_4_data;
  wire [1-1:0] stream_conv2d_24__reduce_reset_data;
  wire [1-1:0] stream_conv2d_24_parameter_6_data;
  wire [32-1:0] stream_conv2d_24_source_7_data;
  wire [1-1:0] stream_conv2d_24_parameter_8_data;
  wire [8-1:0] stream_conv2d_24_source_9_data;
  wire [1-1:0] stream_conv2d_24_parameter_10_data;
  wire [8-1:0] stream_conv2d_24_source_11_data;
  wire [1-1:0] stream_conv2d_24_parameter_12_data;
  wire [8-1:0] stream_conv2d_24_source_13_data;
  wire [1-1:0] stream_conv2d_24_parameter_14_data;
  wire [8-1:0] stream_conv2d_24_source_15_data;
  wire [1-1:0] stream_conv2d_24_parameter_16_data;
  wire [1-1:0] stream_conv2d_24_parameter_17_data;
  wire [5-1:0] stream_conv2d_24_parameter_18_data;
  wire [1-1:0] stream_conv2d_24_parameter_19_data;
  wire [8-1:0] stream_conv2d_24_source_20_data;
  wire [8-1:0] stream_conv2d_24_source_21_data;
  wire [8-1:0] stream_conv2d_24_source_22_data;
  wire [8-1:0] stream_conv2d_24_source_23_data;
  wire [8-1:0] stream_conv2d_24_source_24_data;
  wire [8-1:0] stream_conv2d_24_source_25_data;
  wire [8-1:0] stream_conv2d_24_source_26_data;
  wire [8-1:0] stream_conv2d_24_source_27_data;
  wire [8-1:0] stream_conv2d_24_source_28_data;
  wire [8-1:0] stream_conv2d_24_source_29_data;
  wire [8-1:0] stream_conv2d_24_source_30_data;
  wire [8-1:0] stream_conv2d_24_source_31_data;
  wire [8-1:0] stream_conv2d_24_source_32_data;
  wire [8-1:0] stream_conv2d_24_source_33_data;
  wire [8-1:0] stream_conv2d_24_source_34_data;
  wire [8-1:0] stream_conv2d_24_source_35_data;
  wire [8-1:0] stream_conv2d_24_source_36_data;
  wire [8-1:0] stream_conv2d_24_source_37_data;
  reg __stream_conv2d_24_stream_ivalid_1;
  reg __stream_conv2d_24_stream_ivalid_2;
  reg __stream_conv2d_24_stream_ivalid_3;
  reg __stream_conv2d_24_stream_ivalid_4;
  reg __stream_conv2d_24_stream_ivalid_5;
  reg __stream_conv2d_24_stream_ivalid_6;
  reg __stream_conv2d_24_stream_ivalid_7;
  reg __stream_conv2d_24_stream_ivalid_8;
  reg __stream_conv2d_24_stream_ivalid_9;
  reg __stream_conv2d_24_stream_ivalid_10;
  reg __stream_conv2d_24_stream_ivalid_11;
  reg __stream_conv2d_24_stream_ivalid_12;
  reg __stream_conv2d_24_stream_ivalid_13;
  reg __stream_conv2d_24_stream_ivalid_14;
  reg __stream_conv2d_24_stream_ivalid_15;
  reg __stream_conv2d_24_stream_ivalid_16;
  reg __stream_conv2d_24_stream_ivalid_17;
  reg __stream_conv2d_24_stream_ivalid_18;
  reg __stream_conv2d_24_stream_ivalid_19;
  reg __stream_conv2d_24_stream_ivalid_20;
  reg __stream_conv2d_24_stream_ivalid_21;
  reg __stream_conv2d_24_stream_ivalid_22;
  reg __stream_conv2d_24_stream_ivalid_23;
  reg __stream_conv2d_24_stream_ivalid_24;
  reg __stream_conv2d_24_stream_ivalid_25;
  reg __stream_conv2d_24_stream_ivalid_26;
  reg __stream_conv2d_24_stream_ivalid_27;
  reg __stream_conv2d_24_stream_ivalid_28;
  reg __stream_conv2d_24_stream_ivalid_29;
  reg __stream_conv2d_24_stream_ivalid_30;
  reg __stream_conv2d_24_stream_ivalid_31;
  wire [32-1:0] _slice_data_323;
  assign _slice_data_323 = stream_conv2d_24_source_7_data[6'd31:1'd0];
  wire [32-1:0] _reinterpretcast_src_324;
  assign _reinterpretcast_src_324 = _slice_data_323;
  wire signed [32-1:0] _reinterpretcast_data_324;
  assign _reinterpretcast_data_324 = _reinterpretcast_src_324;
  wire signed [32-1:0] _cond_data_325;
  assign _cond_data_325 = (stream_conv2d_24_parameter_6_data)? _reinterpretcast_data_324 : _reinterpretcast_data_324;
  wire [8-1:0] _slice_data_330;
  assign _slice_data_330 = stream_conv2d_24_source_9_data[4'd7:1'd0];
  wire [8-1:0] _reinterpretcast_src_331;
  assign _reinterpretcast_src_331 = _slice_data_330;
  wire signed [8-1:0] _reinterpretcast_data_331;
  assign _reinterpretcast_data_331 = _reinterpretcast_src_331;
  wire signed [8-1:0] _cond_data_332;
  assign _cond_data_332 = (stream_conv2d_24_parameter_8_data)? _reinterpretcast_data_331 : _reinterpretcast_data_331;
  wire [8-1:0] _slice_data_337;
  assign _slice_data_337 = stream_conv2d_24_source_11_data[4'd7:1'd0];
  wire [8-1:0] _reinterpretcast_src_338;
  assign _reinterpretcast_src_338 = _slice_data_337;
  wire [8-1:0] _reinterpretcast_data_338;
  assign _reinterpretcast_data_338 = _reinterpretcast_src_338;
  wire [8-1:0] _cond_data_339;
  assign _cond_data_339 = (stream_conv2d_24_parameter_10_data)? _reinterpretcast_data_338 : _reinterpretcast_data_338;
  wire [8-1:0] _slice_data_344;
  assign _slice_data_344 = stream_conv2d_24_source_13_data[4'd7:1'd0];
  wire [8-1:0] _reinterpretcast_src_345;
  assign _reinterpretcast_src_345 = _slice_data_344;
  wire [8-1:0] _reinterpretcast_data_345;
  assign _reinterpretcast_data_345 = _reinterpretcast_src_345;
  wire [8-1:0] _cond_data_346;
  assign _cond_data_346 = (stream_conv2d_24_parameter_12_data)? _reinterpretcast_data_345 : _reinterpretcast_data_345;
  wire [8-1:0] _slice_data_351;
  assign _slice_data_351 = stream_conv2d_24_source_15_data[4'd7:1'd0];
  wire [8-1:0] _reinterpretcast_src_352;
  assign _reinterpretcast_src_352 = _slice_data_351;
  wire [8-1:0] _reinterpretcast_data_352;
  assign _reinterpretcast_data_352 = _reinterpretcast_src_352;
  wire [8-1:0] _cond_data_353;
  assign _cond_data_353 = (stream_conv2d_24_parameter_14_data)? _reinterpretcast_data_352 : _reinterpretcast_data_352;
  reg [1-1:0] _eq_data_367;
  reg [1-1:0] _eq_data_371;
  reg [1-1:0] _eq_data_374;
  reg [1-1:0] _eq_data_377;
  reg [1-1:0] _eq_data_381;
  reg [1-1:0] _eq_data_384;
  reg [1-1:0] _eq_data_387;
  reg [1-1:0] _eq_data_391;
  reg [1-1:0] _eq_data_394;
  reg [1-1:0] _eq_data_397;
  reg [1-1:0] _eq_data_401;
  reg [1-1:0] _eq_data_404;
  reg [1-1:0] _eq_data_407;
  reg [1-1:0] _eq_data_411;
  reg [1-1:0] _eq_data_414;
  reg [1-1:0] _eq_data_417;
  reg [1-1:0] _eq_data_421;
  reg [1-1:0] _eq_data_424;
  reg [1-1:0] _eq_data_427;
  reg [1-1:0] _eq_data_431;
  reg [1-1:0] _eq_data_434;
  reg [1-1:0] _eq_data_437;
  reg [1-1:0] _eq_data_441;
  reg [1-1:0] _eq_data_444;
  reg [1-1:0] _eq_data_447;
  reg [1-1:0] _eq_data_451;
  reg [1-1:0] _eq_data_454;
  reg [1-1:0] _eq_data_457;
  reg [1-1:0] _eq_data_461;
  reg [1-1:0] _eq_data_464;
  reg [1-1:0] _eq_data_467;
  reg [1-1:0] _eq_data_471;
  reg [1-1:0] _eq_data_474;
  reg [1-1:0] _eq_data_477;
  reg [1-1:0] _eq_data_481;
  reg [1-1:0] _eq_data_484;
  reg [1-1:0] _eq_data_487;
  reg [1-1:0] _eq_data_491;
  reg [1-1:0] _eq_data_494;
  reg [1-1:0] _eq_data_497;
  reg [1-1:0] _eq_data_501;
  reg [1-1:0] _eq_data_504;
  reg [1-1:0] _eq_data_507;
  reg [1-1:0] _eq_data_511;
  reg [1-1:0] _eq_data_514;
  reg [1-1:0] _eq_data_517;
  reg [1-1:0] _eq_data_521;
  reg [1-1:0] _eq_data_524;
  reg [1-1:0] _eq_data_527;
  reg [1-1:0] _eq_data_531;
  reg [1-1:0] _eq_data_534;
  reg [1-1:0] _eq_data_537;
  reg [1-1:0] _eq_data_541;
  reg [1-1:0] _eq_data_544;
  wire [8-1:0] _reinterpretcast_src_637;
  assign _reinterpretcast_src_637 = stream_conv2d_24_source_29_data;
  wire signed [8-1:0] _reinterpretcast_data_637;
  assign _reinterpretcast_data_637 = _reinterpretcast_src_637;
  wire [8-1:0] _reinterpretcast_src_638;
  assign _reinterpretcast_src_638 = stream_conv2d_24_source_30_data;
  wire signed [8-1:0] _reinterpretcast_data_638;
  assign _reinterpretcast_data_638 = _reinterpretcast_src_638;
  wire [8-1:0] _reinterpretcast_src_639;
  assign _reinterpretcast_src_639 = stream_conv2d_24_source_31_data;
  wire signed [8-1:0] _reinterpretcast_data_639;
  assign _reinterpretcast_data_639 = _reinterpretcast_src_639;
  wire [8-1:0] _reinterpretcast_src_640;
  assign _reinterpretcast_src_640 = stream_conv2d_24_source_32_data;
  wire signed [8-1:0] _reinterpretcast_data_640;
  assign _reinterpretcast_data_640 = _reinterpretcast_src_640;
  wire [8-1:0] _reinterpretcast_src_641;
  assign _reinterpretcast_src_641 = stream_conv2d_24_source_33_data;
  wire signed [8-1:0] _reinterpretcast_data_641;
  assign _reinterpretcast_data_641 = _reinterpretcast_src_641;
  wire [8-1:0] _reinterpretcast_src_642;
  assign _reinterpretcast_src_642 = stream_conv2d_24_source_34_data;
  wire signed [8-1:0] _reinterpretcast_data_642;
  assign _reinterpretcast_data_642 = _reinterpretcast_src_642;
  wire [8-1:0] _reinterpretcast_src_643;
  assign _reinterpretcast_src_643 = stream_conv2d_24_source_35_data;
  wire signed [8-1:0] _reinterpretcast_data_643;
  assign _reinterpretcast_data_643 = _reinterpretcast_src_643;
  wire [8-1:0] _reinterpretcast_src_644;
  assign _reinterpretcast_src_644 = stream_conv2d_24_source_36_data;
  wire signed [8-1:0] _reinterpretcast_data_644;
  assign _reinterpretcast_data_644 = _reinterpretcast_src_644;
  wire [8-1:0] _reinterpretcast_src_645;
  assign _reinterpretcast_src_645 = stream_conv2d_24_source_37_data;
  wire signed [8-1:0] _reinterpretcast_data_645;
  assign _reinterpretcast_data_645 = _reinterpretcast_src_645;
  wire [1-1:0] _pointer_data_646;
  assign _pointer_data_646 = stream_conv2d_24_parameter_3_data[1'sd0];
  wire [1-1:0] _pointer_data_648;
  assign _pointer_data_648 = stream_conv2d_24_parameter_3_data[2'sd1];
  wire [1-1:0] _pointer_data_650;
  assign _pointer_data_650 = stream_conv2d_24_parameter_3_data[3'sd2];
  wire [1-1:0] _pointer_data_652;
  assign _pointer_data_652 = stream_conv2d_24_parameter_3_data[3'sd3];
  wire [1-1:0] _pointer_data_654;
  assign _pointer_data_654 = stream_conv2d_24_parameter_3_data[4'sd4];
  wire [1-1:0] _pointer_data_656;
  assign _pointer_data_656 = stream_conv2d_24_parameter_3_data[4'sd5];
  wire [1-1:0] _pointer_data_658;
  assign _pointer_data_658 = stream_conv2d_24_parameter_3_data[4'sd6];
  wire [1-1:0] _pointer_data_660;
  assign _pointer_data_660 = stream_conv2d_24_parameter_3_data[4'sd7];
  wire [1-1:0] _pointer_data_662;
  assign _pointer_data_662 = stream_conv2d_24_parameter_3_data[5'sd8];
  reg [8-1:0] _plus_data_699;
  reg [8-1:0] _plus_data_718;
  reg [8-1:0] _plus_data_737;
  reg [8-1:0] _plus_data_756;
  reg [8-1:0] _plus_data_775;
  reg [8-1:0] _plus_data_794;
  reg [8-1:0] _plus_data_813;
  reg [8-1:0] _plus_data_832;
  reg [8-1:0] _plus_data_851;
  reg [8-1:0] _plus_data_867;
  reg [8-1:0] _plus_data_886;
  reg [8-1:0] __delay_data_1038__variable_360;
  reg [8-1:0] __delay_data_1039__variable_359;
  reg [8-1:0] __delay_data_1040__variable_358;
  reg [8-1:0] __delay_data_1041__variable_363;
  reg [8-1:0] __delay_data_1042__variable_362;
  reg [8-1:0] __delay_data_1043__variable_361;
  reg [8-1:0] __delay_data_1044__variable_366;
  reg [8-1:0] __delay_data_1045__variable_365;
  reg [8-1:0] __delay_data_1046__variable_364;
  reg [1-1:0] __delay_data_1047_pointer_646;
  reg signed [8-1:0] __delay_data_1048_reinterpretcast_637;
  reg [1-1:0] __delay_data_1049_pointer_648;
  reg signed [8-1:0] __delay_data_1050_reinterpretcast_638;
  reg [1-1:0] __delay_data_1051_pointer_650;
  reg signed [8-1:0] __delay_data_1052_reinterpretcast_639;
  reg [1-1:0] __delay_data_1053_pointer_652;
  reg signed [8-1:0] __delay_data_1054_reinterpretcast_640;
  reg [1-1:0] __delay_data_1055_pointer_654;
  reg signed [8-1:0] __delay_data_1056_reinterpretcast_641;
  reg [1-1:0] __delay_data_1057_pointer_656;
  reg signed [8-1:0] __delay_data_1058_reinterpretcast_642;
  reg [1-1:0] __delay_data_1059_pointer_658;
  reg signed [8-1:0] __delay_data_1060_reinterpretcast_643;
  reg [1-1:0] __delay_data_1061_pointer_660;
  reg signed [8-1:0] __delay_data_1062_reinterpretcast_644;
  reg [1-1:0] __delay_data_1063_pointer_662;
  reg signed [8-1:0] __delay_data_1064_reinterpretcast_645;
  reg [1-1:0] __delay_data_1065__variable_309;
  reg [10-1:0] __delay_data_1090__variable_304;
  reg signed [32-1:0] __delay_data_1103_cond_325;
  reg signed [8-1:0] __delay_data_1122_cond_332;
  wire signed [8-1:0] _cond_data_369;
  assign _cond_data_369 = (_eq_data_367)? __delay_data_1038__variable_360 : 1'sd0;
  wire signed [8-1:0] _cond_data_373;
  assign _cond_data_373 = (_eq_data_371)? __delay_data_1039__variable_359 : _cond_data_369;
  wire signed [8-1:0] _cond_data_376;
  assign _cond_data_376 = (_eq_data_374)? __delay_data_1040__variable_358 : _cond_data_373;
  wire signed [8-1:0] _cond_data_379;
  assign _cond_data_379 = (_eq_data_377)? __delay_data_1040__variable_358 : 1'sd0;
  wire signed [8-1:0] _cond_data_383;
  assign _cond_data_383 = (_eq_data_381)? __delay_data_1038__variable_360 : _cond_data_379;
  wire signed [8-1:0] _cond_data_386;
  assign _cond_data_386 = (_eq_data_384)? __delay_data_1039__variable_359 : _cond_data_383;
  wire signed [8-1:0] _cond_data_389;
  assign _cond_data_389 = (_eq_data_387)? __delay_data_1039__variable_359 : 1'sd0;
  wire signed [8-1:0] _cond_data_393;
  assign _cond_data_393 = (_eq_data_391)? __delay_data_1040__variable_358 : _cond_data_389;
  wire signed [8-1:0] _cond_data_396;
  assign _cond_data_396 = (_eq_data_394)? __delay_data_1038__variable_360 : _cond_data_393;
  wire signed [8-1:0] _cond_data_399;
  assign _cond_data_399 = (_eq_data_397)? __delay_data_1041__variable_363 : 1'sd0;
  wire signed [8-1:0] _cond_data_403;
  assign _cond_data_403 = (_eq_data_401)? __delay_data_1042__variable_362 : _cond_data_399;
  wire signed [8-1:0] _cond_data_406;
  assign _cond_data_406 = (_eq_data_404)? __delay_data_1043__variable_361 : _cond_data_403;
  wire signed [8-1:0] _cond_data_409;
  assign _cond_data_409 = (_eq_data_407)? __delay_data_1043__variable_361 : 1'sd0;
  wire signed [8-1:0] _cond_data_413;
  assign _cond_data_413 = (_eq_data_411)? __delay_data_1041__variable_363 : _cond_data_409;
  wire signed [8-1:0] _cond_data_416;
  assign _cond_data_416 = (_eq_data_414)? __delay_data_1042__variable_362 : _cond_data_413;
  wire signed [8-1:0] _cond_data_419;
  assign _cond_data_419 = (_eq_data_417)? __delay_data_1042__variable_362 : 1'sd0;
  wire signed [8-1:0] _cond_data_423;
  assign _cond_data_423 = (_eq_data_421)? __delay_data_1043__variable_361 : _cond_data_419;
  wire signed [8-1:0] _cond_data_426;
  assign _cond_data_426 = (_eq_data_424)? __delay_data_1041__variable_363 : _cond_data_423;
  wire signed [8-1:0] _cond_data_429;
  assign _cond_data_429 = (_eq_data_427)? __delay_data_1044__variable_366 : 1'sd0;
  wire signed [8-1:0] _cond_data_433;
  assign _cond_data_433 = (_eq_data_431)? __delay_data_1045__variable_365 : _cond_data_429;
  wire signed [8-1:0] _cond_data_436;
  assign _cond_data_436 = (_eq_data_434)? __delay_data_1046__variable_364 : _cond_data_433;
  wire signed [8-1:0] _cond_data_439;
  assign _cond_data_439 = (_eq_data_437)? __delay_data_1046__variable_364 : 1'sd0;
  wire signed [8-1:0] _cond_data_443;
  assign _cond_data_443 = (_eq_data_441)? __delay_data_1044__variable_366 : _cond_data_439;
  wire signed [8-1:0] _cond_data_446;
  assign _cond_data_446 = (_eq_data_444)? __delay_data_1045__variable_365 : _cond_data_443;
  wire signed [8-1:0] _cond_data_449;
  assign _cond_data_449 = (_eq_data_447)? __delay_data_1045__variable_365 : 1'sd0;
  wire signed [8-1:0] _cond_data_453;
  assign _cond_data_453 = (_eq_data_451)? __delay_data_1046__variable_364 : _cond_data_449;
  wire signed [8-1:0] _cond_data_456;
  assign _cond_data_456 = (_eq_data_454)? __delay_data_1044__variable_366 : _cond_data_453;
  wire signed [8-1:0] _cond_data_459;
  assign _cond_data_459 = (_eq_data_457)? _cond_data_436 : 1'sd0;
  wire signed [8-1:0] _cond_data_463;
  assign _cond_data_463 = (_eq_data_461)? _cond_data_406 : _cond_data_459;
  wire signed [8-1:0] _cond_data_466;
  assign _cond_data_466 = (_eq_data_464)? _cond_data_376 : _cond_data_463;
  wire signed [8-1:0] _cond_data_469;
  assign _cond_data_469 = (_eq_data_467)? _cond_data_376 : 1'sd0;
  wire signed [8-1:0] _cond_data_473;
  assign _cond_data_473 = (_eq_data_471)? _cond_data_436 : _cond_data_469;
  wire signed [8-1:0] _cond_data_476;
  assign _cond_data_476 = (_eq_data_474)? _cond_data_406 : _cond_data_473;
  wire signed [8-1:0] _cond_data_479;
  assign _cond_data_479 = (_eq_data_477)? _cond_data_406 : 1'sd0;
  wire signed [8-1:0] _cond_data_483;
  assign _cond_data_483 = (_eq_data_481)? _cond_data_376 : _cond_data_479;
  wire signed [8-1:0] _cond_data_486;
  assign _cond_data_486 = (_eq_data_484)? _cond_data_436 : _cond_data_483;
  wire signed [8-1:0] _cond_data_489;
  assign _cond_data_489 = (_eq_data_487)? _cond_data_446 : 1'sd0;
  wire signed [8-1:0] _cond_data_493;
  assign _cond_data_493 = (_eq_data_491)? _cond_data_416 : _cond_data_489;
  wire signed [8-1:0] _cond_data_496;
  assign _cond_data_496 = (_eq_data_494)? _cond_data_386 : _cond_data_493;
  wire signed [8-1:0] _cond_data_499;
  assign _cond_data_499 = (_eq_data_497)? _cond_data_386 : 1'sd0;
  wire signed [8-1:0] _cond_data_503;
  assign _cond_data_503 = (_eq_data_501)? _cond_data_446 : _cond_data_499;
  wire signed [8-1:0] _cond_data_506;
  assign _cond_data_506 = (_eq_data_504)? _cond_data_416 : _cond_data_503;
  wire signed [8-1:0] _cond_data_509;
  assign _cond_data_509 = (_eq_data_507)? _cond_data_416 : 1'sd0;
  wire signed [8-1:0] _cond_data_513;
  assign _cond_data_513 = (_eq_data_511)? _cond_data_386 : _cond_data_509;
  wire signed [8-1:0] _cond_data_516;
  assign _cond_data_516 = (_eq_data_514)? _cond_data_446 : _cond_data_513;
  wire signed [8-1:0] _cond_data_519;
  assign _cond_data_519 = (_eq_data_517)? _cond_data_456 : 1'sd0;
  wire signed [8-1:0] _cond_data_523;
  assign _cond_data_523 = (_eq_data_521)? _cond_data_426 : _cond_data_519;
  wire signed [8-1:0] _cond_data_526;
  assign _cond_data_526 = (_eq_data_524)? _cond_data_396 : _cond_data_523;
  wire signed [8-1:0] _cond_data_529;
  assign _cond_data_529 = (_eq_data_527)? _cond_data_396 : 1'sd0;
  wire signed [8-1:0] _cond_data_533;
  assign _cond_data_533 = (_eq_data_531)? _cond_data_456 : _cond_data_529;
  wire signed [8-1:0] _cond_data_536;
  assign _cond_data_536 = (_eq_data_534)? _cond_data_426 : _cond_data_533;
  wire signed [8-1:0] _cond_data_539;
  assign _cond_data_539 = (_eq_data_537)? _cond_data_426 : 1'sd0;
  wire signed [8-1:0] _cond_data_543;
  assign _cond_data_543 = (_eq_data_541)? _cond_data_396 : _cond_data_539;
  wire signed [8-1:0] _cond_data_546;
  assign _cond_data_546 = (_eq_data_544)? _cond_data_456 : _cond_data_543;
  wire signed [8-1:0] _reinterpretcast_src_583;
  assign _reinterpretcast_src_583 = _cond_data_466;
  wire signed [8-1:0] _reinterpretcast_data_583;
  assign _reinterpretcast_data_583 = _reinterpretcast_src_583;
  wire signed [8-1:0] _reinterpretcast_src_584;
  assign _reinterpretcast_src_584 = _cond_data_496;
  wire signed [8-1:0] _reinterpretcast_data_584;
  assign _reinterpretcast_data_584 = _reinterpretcast_src_584;
  wire signed [8-1:0] _reinterpretcast_src_585;
  assign _reinterpretcast_src_585 = _cond_data_526;
  wire signed [8-1:0] _reinterpretcast_data_585;
  assign _reinterpretcast_data_585 = _reinterpretcast_src_585;
  wire signed [8-1:0] _reinterpretcast_src_586;
  assign _reinterpretcast_src_586 = _cond_data_476;
  wire signed [8-1:0] _reinterpretcast_data_586;
  assign _reinterpretcast_data_586 = _reinterpretcast_src_586;
  wire signed [8-1:0] _reinterpretcast_src_587;
  assign _reinterpretcast_src_587 = _cond_data_506;
  wire signed [8-1:0] _reinterpretcast_data_587;
  assign _reinterpretcast_data_587 = _reinterpretcast_src_587;
  wire signed [8-1:0] _reinterpretcast_src_588;
  assign _reinterpretcast_src_588 = _cond_data_536;
  wire signed [8-1:0] _reinterpretcast_data_588;
  assign _reinterpretcast_data_588 = _reinterpretcast_src_588;
  wire signed [8-1:0] _reinterpretcast_src_589;
  assign _reinterpretcast_src_589 = _cond_data_486;
  wire signed [8-1:0] _reinterpretcast_data_589;
  assign _reinterpretcast_data_589 = _reinterpretcast_src_589;
  wire signed [8-1:0] _reinterpretcast_src_590;
  assign _reinterpretcast_src_590 = _cond_data_516;
  wire signed [8-1:0] _reinterpretcast_data_590;
  assign _reinterpretcast_data_590 = _reinterpretcast_src_590;
  wire signed [8-1:0] _reinterpretcast_src_591;
  assign _reinterpretcast_src_591 = _cond_data_546;
  wire signed [8-1:0] _reinterpretcast_data_591;
  assign _reinterpretcast_data_591 = _reinterpretcast_src_591;
  wire signed [8-1:0] _cond_data_665;
  assign _cond_data_665 = (__delay_data_1047_pointer_646)? 1'sd0 : _reinterpretcast_data_583;
  wire signed [8-1:0] _cond_data_667;
  assign _cond_data_667 = (__delay_data_1049_pointer_648)? 1'sd0 : _reinterpretcast_data_584;
  wire signed [8-1:0] _cond_data_669;
  assign _cond_data_669 = (__delay_data_1051_pointer_650)? 1'sd0 : _reinterpretcast_data_585;
  wire signed [8-1:0] _cond_data_671;
  assign _cond_data_671 = (__delay_data_1053_pointer_652)? 1'sd0 : _reinterpretcast_data_586;
  wire signed [8-1:0] _cond_data_673;
  assign _cond_data_673 = (__delay_data_1055_pointer_654)? 1'sd0 : _reinterpretcast_data_587;
  wire signed [8-1:0] _cond_data_675;
  assign _cond_data_675 = (__delay_data_1057_pointer_656)? 1'sd0 : _reinterpretcast_data_588;
  wire signed [8-1:0] _cond_data_677;
  assign _cond_data_677 = (__delay_data_1059_pointer_658)? 1'sd0 : _reinterpretcast_data_589;
  wire signed [8-1:0] _cond_data_679;
  assign _cond_data_679 = (__delay_data_1061_pointer_660)? 1'sd0 : _reinterpretcast_data_590;
  wire signed [8-1:0] _cond_data_681;
  assign _cond_data_681 = (__delay_data_1063_pointer_662)? 1'sd0 : _reinterpretcast_data_591;
  reg signed [8-1:0] __variable_wdata_108;
  assign mul_5_x_data = __variable_wdata_108;
  reg signed [8-1:0] __variable_wdata_109;
  assign mul_5_y_data = __variable_wdata_109;
  reg [4-1:0] __variable_wdata_110;
  assign mul_5_rshift_data = __variable_wdata_110;
  reg signed [8-1:0] __variable_wdata_129;
  assign mul_6_x_data = __variable_wdata_129;
  reg signed [8-1:0] __variable_wdata_130;
  assign mul_6_y_data = __variable_wdata_130;
  reg [4-1:0] __variable_wdata_131;
  assign mul_6_rshift_data = __variable_wdata_131;
  assign _mul_6_is_root = ((_stream_conv2d_24_busy)? 0 : 1) && 1;
  assign _mul_6_stream_oready = ((_stream_conv2d_24_busy)? _stream_conv2d_24_stream_oready : 1) && _mul_6_stream_internal_oready;
  reg signed [8-1:0] __variable_wdata_150;
  assign mul_7_x_data = __variable_wdata_150;
  reg signed [8-1:0] __variable_wdata_151;
  assign mul_7_y_data = __variable_wdata_151;
  reg [4-1:0] __variable_wdata_152;
  assign mul_7_rshift_data = __variable_wdata_152;
  assign _mul_7_is_root = ((_stream_conv2d_24_busy)? 0 : 1) && 1;
  assign _mul_7_stream_oready = ((_stream_conv2d_24_busy)? _stream_conv2d_24_stream_oready : 1) && _mul_7_stream_internal_oready;
  reg signed [8-1:0] __variable_wdata_171;
  assign mul_8_x_data = __variable_wdata_171;
  reg signed [8-1:0] __variable_wdata_172;
  assign mul_8_y_data = __variable_wdata_172;
  reg [4-1:0] __variable_wdata_173;
  assign mul_8_rshift_data = __variable_wdata_173;
  assign _mul_8_is_root = ((_stream_conv2d_24_busy)? 0 : 1) && 1;
  assign _mul_8_stream_oready = ((_stream_conv2d_24_busy)? _stream_conv2d_24_stream_oready : 1) && _mul_8_stream_internal_oready;
  reg signed [8-1:0] __variable_wdata_192;
  assign mul_9_x_data = __variable_wdata_192;
  reg signed [8-1:0] __variable_wdata_193;
  assign mul_9_y_data = __variable_wdata_193;
  reg [4-1:0] __variable_wdata_194;
  assign mul_9_rshift_data = __variable_wdata_194;
  assign _mul_9_is_root = ((_stream_conv2d_24_busy)? 0 : 1) && 1;
  assign _mul_9_stream_oready = ((_stream_conv2d_24_busy)? _stream_conv2d_24_stream_oready : 1) && _mul_9_stream_internal_oready;
  reg signed [8-1:0] __variable_wdata_213;
  assign mul_10_x_data = __variable_wdata_213;
  reg signed [8-1:0] __variable_wdata_214;
  assign mul_10_y_data = __variable_wdata_214;
  reg [4-1:0] __variable_wdata_215;
  assign mul_10_rshift_data = __variable_wdata_215;
  assign _mul_10_is_root = ((_stream_conv2d_24_busy)? 0 : 1) && 1;
  assign _mul_10_stream_oready = ((_stream_conv2d_24_busy)? _stream_conv2d_24_stream_oready : 1) && _mul_10_stream_internal_oready;
  reg signed [8-1:0] __variable_wdata_234;
  assign mul_11_x_data = __variable_wdata_234;
  reg signed [8-1:0] __variable_wdata_235;
  assign mul_11_y_data = __variable_wdata_235;
  reg [4-1:0] __variable_wdata_236;
  assign mul_11_rshift_data = __variable_wdata_236;
  assign _mul_11_is_root = ((_stream_conv2d_24_busy)? 0 : 1) && 1;
  assign _mul_11_stream_oready = ((_stream_conv2d_24_busy)? _stream_conv2d_24_stream_oready : 1) && _mul_11_stream_internal_oready;
  reg signed [8-1:0] __variable_wdata_255;
  assign mul_12_x_data = __variable_wdata_255;
  reg signed [8-1:0] __variable_wdata_256;
  assign mul_12_y_data = __variable_wdata_256;
  reg [4-1:0] __variable_wdata_257;
  assign mul_12_rshift_data = __variable_wdata_257;
  assign _mul_12_is_root = ((_stream_conv2d_24_busy)? 0 : 1) && 1;
  assign _mul_12_stream_oready = ((_stream_conv2d_24_busy)? _stream_conv2d_24_stream_oready : 1) && _mul_12_stream_internal_oready;
  reg signed [8-1:0] __variable_wdata_276;
  assign mul_13_x_data = __variable_wdata_276;
  reg signed [8-1:0] __variable_wdata_277;
  assign mul_13_y_data = __variable_wdata_277;
  reg [4-1:0] __variable_wdata_278;
  assign mul_13_rshift_data = __variable_wdata_278;
  assign _mul_13_is_root = ((_stream_conv2d_24_busy)? 0 : 1) && 1;
  assign _mul_13_stream_oready = ((_stream_conv2d_24_busy)? _stream_conv2d_24_stream_oready : 1) && _mul_13_stream_internal_oready;
  reg [1-1:0] __delay_data_1066__delay_1065__variable_309;
  reg [8-1:0] __delay_data_1078_plus_867;
  reg [10-1:0] __delay_data_1091__delay_1090__variable_304;
  reg signed [32-1:0] __delay_data_1104__delay_1103_cond_325;
  reg signed [8-1:0] __delay_data_1123__delay_1122_cond_332;
  reg [8-1:0] __delay_data_1142_plus_886;
  reg [1-1:0] __delay_data_1067__delay_1066__delay_1065__variable_309;
  reg [8-1:0] __delay_data_1079__delay_1078_plus_867;
  reg [10-1:0] __delay_data_1092__delay_1091__delay_1090__variable_304;
  reg signed [32-1:0] __delay_data_1105__delay_1104__delay_1103_cond_325;
  reg signed [8-1:0] __delay_data_1124__delay_1123__delay_1122_cond_332;
  reg [8-1:0] __delay_data_1143__delay_1142_plus_886;
  reg [1-1:0] __delay_data_1068__delay_1067__delay_1066____variable_309;
  reg [8-1:0] __delay_data_1080__delay_1079__delay_1078_plus_867;
  reg [10-1:0] __delay_data_1093__delay_1092__delay_1091____variable_304;
  reg signed [32-1:0] __delay_data_1106__delay_1105__delay_1104__delay_1103_cond_325;
  reg signed [8-1:0] __delay_data_1125__delay_1124__delay_1123__delay_1122_cond_332;
  reg [8-1:0] __delay_data_1144__delay_1143__delay_1142_plus_886;
  reg [1-1:0] __delay_data_1069__delay_1068__delay_1067____variable_309;
  reg [8-1:0] __delay_data_1081__delay_1080__delay_1079__delay_1078_plus_867;
  reg [10-1:0] __delay_data_1094__delay_1093__delay_1092____variable_304;
  reg signed [32-1:0] __delay_data_1107__delay_1106__delay_1105__delay_1104___cond_325;
  reg signed [8-1:0] __delay_data_1126__delay_1125__delay_1124__delay_1123___cond_332;
  reg [8-1:0] __delay_data_1145__delay_1144__delay_1143__delay_1142_plus_886;
  reg [1-1:0] __delay_data_1070__delay_1069__delay_1068____variable_309;
  reg [8-1:0] __delay_data_1082__delay_1081__delay_1080__delay_1079___plus_867;
  reg [10-1:0] __delay_data_1095__delay_1094__delay_1093____variable_304;
  reg signed [32-1:0] __delay_data_1108__delay_1107__delay_1106__delay_1105___cond_325;
  reg signed [8-1:0] __delay_data_1127__delay_1126__delay_1125__delay_1124___cond_332;
  reg [8-1:0] __delay_data_1146__delay_1145__delay_1144__delay_1143___plus_886;
  reg [1-1:0] __delay_data_1071__delay_1070__delay_1069____variable_309;
  reg [8-1:0] __delay_data_1083__delay_1082__delay_1081__delay_1080___plus_867;
  reg [10-1:0] __delay_data_1096__delay_1095__delay_1094____variable_304;
  reg signed [32-1:0] __delay_data_1109__delay_1108__delay_1107__delay_1106___cond_325;
  reg signed [8-1:0] __delay_data_1128__delay_1127__delay_1126__delay_1125___cond_332;
  reg [8-1:0] __delay_data_1147__delay_1146__delay_1145__delay_1144___plus_886;
  reg [1-1:0] __delay_data_1072__delay_1071__delay_1070____variable_309;
  reg [8-1:0] __delay_data_1084__delay_1083__delay_1082__delay_1081___plus_867;
  reg [10-1:0] __delay_data_1097__delay_1096__delay_1095____variable_304;
  reg signed [32-1:0] __delay_data_1110__delay_1109__delay_1108__delay_1107___cond_325;
  reg signed [8-1:0] __delay_data_1129__delay_1128__delay_1127__delay_1126___cond_332;
  reg [8-1:0] __delay_data_1148__delay_1147__delay_1146__delay_1145___plus_886;
  reg [1-1:0] __delay_data_1073__delay_1072__delay_1071____variable_309;
  reg [8-1:0] __delay_data_1085__delay_1084__delay_1083__delay_1082___plus_867;
  reg [10-1:0] __delay_data_1098__delay_1097__delay_1096____variable_304;
  reg signed [32-1:0] __delay_data_1111__delay_1110__delay_1109__delay_1108___cond_325;
  reg signed [8-1:0] __delay_data_1130__delay_1129__delay_1128__delay_1127___cond_332;
  reg [8-1:0] __delay_data_1149__delay_1148__delay_1147__delay_1146___plus_886;
  reg [1-1:0] __delay_data_1074__delay_1073__delay_1072____variable_309;
  reg [8-1:0] __delay_data_1086__delay_1085__delay_1084__delay_1083___plus_867;
  reg [10-1:0] __delay_data_1099__delay_1098__delay_1097____variable_304;
  reg signed [32-1:0] __delay_data_1112__delay_1111__delay_1110__delay_1109___cond_325;
  reg signed [8-1:0] __delay_data_1131__delay_1130__delay_1129__delay_1128___cond_332;
  reg [8-1:0] __delay_data_1150__delay_1149__delay_1148__delay_1147___plus_886;
  wire signed [16-1:0] __substreamoutput_data_700;
  assign __substreamoutput_data_700 = mul_5_z_data;
  wire signed [16-1:0] __substreamoutput_data_719;
  assign __substreamoutput_data_719 = mul_6_z_data;
  wire signed [16-1:0] __substreamoutput_data_738;
  assign __substreamoutput_data_738 = mul_7_z_data;
  wire signed [16-1:0] __substreamoutput_data_757;
  assign __substreamoutput_data_757 = mul_8_z_data;
  wire signed [16-1:0] __substreamoutput_data_776;
  assign __substreamoutput_data_776 = mul_9_z_data;
  wire signed [16-1:0] __substreamoutput_data_795;
  assign __substreamoutput_data_795 = mul_10_z_data;
  wire signed [16-1:0] __substreamoutput_data_814;
  assign __substreamoutput_data_814 = mul_11_z_data;
  wire signed [16-1:0] __substreamoutput_data_833;
  assign __substreamoutput_data_833 = mul_12_z_data;
  wire signed [16-1:0] __substreamoutput_data_852;
  assign __substreamoutput_data_852 = mul_13_z_data;
  reg signed [32-1:0] __variable_wdata_60;
  assign add_tree_3_var0_data = __variable_wdata_60;
  reg signed [32-1:0] __variable_wdata_61;
  assign add_tree_3_var1_data = __variable_wdata_61;
  reg signed [32-1:0] __variable_wdata_62;
  assign add_tree_3_var2_data = __variable_wdata_62;
  reg signed [32-1:0] __variable_wdata_63;
  assign add_tree_3_var3_data = __variable_wdata_63;
  reg signed [32-1:0] __variable_wdata_64;
  assign add_tree_3_var4_data = __variable_wdata_64;
  reg signed [32-1:0] __variable_wdata_65;
  assign add_tree_3_var5_data = __variable_wdata_65;
  reg signed [32-1:0] __variable_wdata_66;
  assign add_tree_3_var6_data = __variable_wdata_66;
  reg signed [32-1:0] __variable_wdata_67;
  assign add_tree_3_var7_data = __variable_wdata_67;
  reg signed [32-1:0] __variable_wdata_68;
  assign add_tree_3_var8_data = __variable_wdata_68;
  assign _add_tree_3_is_root = ((_stream_conv2d_24_busy)? 0 : 1) && 1;
  assign _add_tree_3_stream_oready = ((_stream_conv2d_24_busy)? _stream_conv2d_24_stream_oready : 1) && _add_tree_3_stream_internal_oready;
  reg [1-1:0] __delay_data_1075__delay_1074__delay_1073____variable_309;
  reg [8-1:0] __delay_data_1087__delay_1086__delay_1085__delay_1084___plus_867;
  reg [10-1:0] __delay_data_1100__delay_1099__delay_1098____variable_304;
  reg signed [32-1:0] __delay_data_1113__delay_1112__delay_1111__delay_1110___cond_325;
  reg signed [8-1:0] __delay_data_1132__delay_1131__delay_1130__delay_1129___cond_332;
  reg [8-1:0] __delay_data_1151__delay_1150__delay_1149__delay_1148___plus_886;
  reg [1-1:0] __delay_data_1076__delay_1075__delay_1074____variable_309;
  reg [8-1:0] __delay_data_1088__delay_1087__delay_1086__delay_1085___plus_867;
  reg [10-1:0] __delay_data_1101__delay_1100__delay_1099____variable_304;
  reg signed [32-1:0] __delay_data_1114__delay_1113__delay_1112__delay_1111___cond_325;
  reg signed [8-1:0] __delay_data_1133__delay_1132__delay_1131__delay_1130___cond_332;
  reg [8-1:0] __delay_data_1152__delay_1151__delay_1150__delay_1149___plus_886;
  reg [1-1:0] __delay_data_1077__delay_1076__delay_1075____variable_309;
  reg [8-1:0] __delay_data_1089__delay_1088__delay_1087__delay_1086___plus_867;
  reg [10-1:0] __delay_data_1102__delay_1101__delay_1100____variable_304;
  reg signed [32-1:0] __delay_data_1115__delay_1114__delay_1113__delay_1112___cond_325;
  reg signed [8-1:0] __delay_data_1134__delay_1133__delay_1132__delay_1131___cond_332;
  reg [8-1:0] __delay_data_1153__delay_1152__delay_1151__delay_1150___plus_886;
  wire signed [32-1:0] __substreamoutput_data_854;
  assign __substreamoutput_data_854 = add_tree_3_sum_data;
  reg [1-1:0] __variable_wdata_51;
  assign acc_1__reduce_reset_data = __variable_wdata_51;
  reg signed [32-1:0] __variable_wdata_36;
  assign acc_1_x_data = __variable_wdata_36;
  reg [6-1:0] __variable_wdata_37;
  assign acc_1_rshift_data = __variable_wdata_37;
  reg [32-1:0] __variable_wdata_38;
  assign acc_1_size_data = __variable_wdata_38;
  reg signed [32-1:0] __delay_data_1116__delay_1115__delay_1114__delay_1113___cond_325;
  reg signed [8-1:0] __delay_data_1135__delay_1134__delay_1133__delay_1132___cond_332;
  reg [8-1:0] __delay_data_1154__delay_1153__delay_1152__delay_1151___plus_886;
  reg signed [32-1:0] __delay_data_1117__delay_1116__delay_1115__delay_1114___cond_325;
  reg signed [8-1:0] __delay_data_1136__delay_1135__delay_1134__delay_1133___cond_332;
  reg [8-1:0] __delay_data_1155__delay_1154__delay_1153__delay_1152___plus_886;
  reg signed [32-1:0] __delay_data_1118__delay_1117__delay_1116__delay_1115___cond_325;
  reg signed [8-1:0] __delay_data_1137__delay_1136__delay_1135__delay_1134___cond_332;
  reg [8-1:0] __delay_data_1156__delay_1155__delay_1154__delay_1153___plus_886;
  reg signed [32-1:0] __delay_data_1119__delay_1118__delay_1117__delay_1116___cond_325;
  reg signed [8-1:0] __delay_data_1138__delay_1137__delay_1136__delay_1135___cond_332;
  reg [8-1:0] __delay_data_1157__delay_1156__delay_1155__delay_1154___plus_886;
  reg signed [32-1:0] __delay_data_1120__delay_1119__delay_1118__delay_1117___cond_325;
  reg signed [8-1:0] __delay_data_1139__delay_1138__delay_1137__delay_1136___cond_332;
  reg [8-1:0] __delay_data_1158__delay_1157__delay_1156__delay_1155___plus_886;
  reg signed [32-1:0] __delay_data_1121__delay_1120__delay_1119__delay_1118___cond_325;
  reg signed [8-1:0] __delay_data_1140__delay_1139__delay_1138__delay_1137___cond_332;
  reg [8-1:0] __delay_data_1159__delay_1158__delay_1157__delay_1156___plus_886;
  wire signed [32-1:0] __substreamoutput_data_868;
  assign __substreamoutput_data_868 = acc_1_sum_data;
  wire [1-1:0] __substreamoutput_data_869;
  assign __substreamoutput_data_869 = acc_1_valid_data;
  reg signed [32-1:0] _plus_data_870;
  reg signed [8-1:0] __delay_data_1141__delay_1140__delay_1139__delay_1138___cond_332;
  reg [8-1:0] __delay_data_1160__delay_1159__delay_1158__delay_1157___plus_886;
  reg [1-1:0] __delay_data_1162__substreamoutput_869;
  reg signed [32-1:0] __variable_wdata_74;
  assign mul_rshift_round_clip_4_x_data = __variable_wdata_74;
  reg signed [8-1:0] __variable_wdata_75;
  assign mul_rshift_round_clip_4_y_data = __variable_wdata_75;
  reg [6-1:0] __variable_wdata_76;
  assign mul_rshift_round_clip_4_rshift_data = __variable_wdata_76;
  assign _stream_conv2d_24_stream_internal_oready = ((_stream_conv2d_24_busy)? _mul_rshift_round_clip_4_stream_internal_oready : 1) && (((_stream_conv2d_24_busy)? _acc_1_stream_internal_oready : 1) && (((_stream_conv2d_24_busy)? _add_tree_3_stream_internal_oready : 1) && (((_stream_conv2d_24_busy)? _mul_13_stream_internal_oready : 1) && (((_stream_conv2d_24_busy)? _mul_12_stream_internal_oready : 1) && (((_stream_conv2d_24_busy)? _mul_11_stream_internal_oready : 1) && (((_stream_conv2d_24_busy)? _mul_10_stream_internal_oready : 1) && (((_stream_conv2d_24_busy)? _mul_9_stream_internal_oready : 1) && (((_stream_conv2d_24_busy)? _mul_8_stream_internal_oready : 1) && (((_stream_conv2d_24_busy)? _mul_7_stream_internal_oready : 1) && (((_stream_conv2d_24_busy)? _mul_6_stream_internal_oready : 1) && (((_stream_conv2d_24_busy)? _mul_5_stream_internal_oready : 1) && 1)))))))))));
  reg [1-1:0] __delay_data_1163__delay_1162__substreamoutput_869;
  reg [1-1:0] __delay_data_1164__delay_1163__delay_1162__substreamoutput_869;
  reg [1-1:0] __delay_data_1165__delay_1164__delay_1163____substreamoutput_869;
  reg [1-1:0] __delay_data_1166__delay_1165__delay_1164____substreamoutput_869;
  reg [1-1:0] __delay_data_1167__delay_1166__delay_1165____substreamoutput_869;
  reg [1-1:0] __delay_data_1168__delay_1167__delay_1166____substreamoutput_869;
  reg [1-1:0] __delay_data_1169__delay_1168__delay_1167____substreamoutput_869;
  reg [1-1:0] __delay_data_1170__delay_1169__delay_1168____substreamoutput_869;
  reg [1-1:0] __delay_data_1171__delay_1170__delay_1169____substreamoutput_869;
  wire signed [8-1:0] __substreamoutput_data_887;
  assign __substreamoutput_data_887 = mul_rshift_round_clip_4_z_data;
  reg [1-1:0] _greaterthan_data_889;
  reg signed [8-1:0] __delay_data_1161__substreamoutput_887;
  reg [1-1:0] __delay_data_1172__delay_1171__delay_1170____substreamoutput_869;
  reg signed [8-1:0] _cond_data_891;
  reg [1-1:0] __delay_data_1173__delay_1172__delay_1171____substreamoutput_869;
  wire signed [8-1:0] _reinterpretcast_src_892;
  assign _reinterpretcast_src_892 = _cond_data_891;
  wire signed [8-1:0] _reinterpretcast_data_892;
  assign _reinterpretcast_data_892 = _reinterpretcast_src_892;
  wire signed [8-1:0] stream_conv2d_24_sink_50_data;
  assign stream_conv2d_24_sink_50_data = _reinterpretcast_data_892;
  wire [1-1:0] stream_conv2d_24_sink_51_data;
  assign stream_conv2d_24_sink_51_data = __delay_data_1173__delay_1172__delay_1171____substreamoutput_869;
  wire _set_flag_397;
  assign _set_flag_397 = conv2d_24_comp_fsm == 3;
  reg [10-1:0] __variable_wdata_304;
  assign stream_conv2d_24_parameter_0_data = __variable_wdata_304;
  wire _set_flag_398;
  assign _set_flag_398 = conv2d_24_comp_fsm == 3;
  reg [2-1:0] __variable_wdata_305;
  assign stream_conv2d_24_parameter_1_data = __variable_wdata_305;
  wire _set_flag_399;
  assign _set_flag_399 = conv2d_24_comp_fsm == 3;
  reg [2-1:0] __variable_wdata_306;
  assign stream_conv2d_24_parameter_2_data = __variable_wdata_306;
  wire _set_flag_400;
  assign _set_flag_400 = conv2d_24_comp_fsm == 3;
  reg [9-1:0] __variable_wdata_307;
  assign stream_conv2d_24_parameter_3_data = __variable_wdata_307;
  wire _set_flag_401;
  assign _set_flag_401 = conv2d_24_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_308;
  assign stream_conv2d_24_parameter_4_data = __variable_wdata_308;
  wire _set_flag_402;
  assign _set_flag_402 = conv2d_24_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_319;
  assign stream_conv2d_24_parameter_6_data = __variable_wdata_319;
  reg [32-1:0] _source_stream_conv2d_24_source_7_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_24_source_7_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_24_source_7_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_24_source_7_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_24_source_7_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_24_source_7_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_24_source_7_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_24_source_7_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_24_source_7_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_24_source_7_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_24_source_7_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_24_source_7_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_24_source_7_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_24_source_7_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_24_source_7_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_24_source_7_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_24_source_7_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_24_source_7_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_24_source_7_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_24_source_7_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_24_source_7_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_24_source_7_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_24_source_7_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_24_source_7_pat_stride_buf_3;
  wire _set_flag_403;
  assign _set_flag_403 = conv2d_24_comp_fsm == 3;
  localparam _tmp_404 = 1;
  wire [_tmp_404-1:0] _tmp_405;
  assign _tmp_405 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_7_source_ram_renable && (_stream_conv2d_24_source_7_source_sel == 1);
  reg [_tmp_404-1:0] __tmp_405_1;
  assign _stream_conv2d_24_source_7_source_ram_rdata = (_stream_conv2d_24_source_7_source_sel == 1)? ram_w32_l4096_id0_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_320;
  assign stream_conv2d_24_source_7_data = __variable_wdata_320;
  reg [32-1:0] _stream_conv2d_24_source_7_source_pat_fsm_0;
  localparam _stream_conv2d_24_source_7_source_pat_fsm_0_init = 0;
  wire [32-1:0] _stream_conv2d_24_source_7_source_pat_all_offset;
  assign _stream_conv2d_24_source_7_source_pat_all_offset = _stream_conv2d_24_source_7_source_offset_buf + _source_stream_conv2d_24_source_7_pat_cur_offset_0 + _source_stream_conv2d_24_source_7_pat_cur_offset_1 + _source_stream_conv2d_24_source_7_pat_cur_offset_2 + _source_stream_conv2d_24_source_7_pat_cur_offset_3;
  wire _set_flag_406;
  assign _set_flag_406 = conv2d_24_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_326;
  assign stream_conv2d_24_parameter_8_data = __variable_wdata_326;
  reg [32-1:0] _source_stream_conv2d_24_source_9_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_24_source_9_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_24_source_9_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_24_source_9_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_24_source_9_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_24_source_9_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_24_source_9_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_24_source_9_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_24_source_9_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_24_source_9_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_24_source_9_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_24_source_9_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_24_source_9_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_24_source_9_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_24_source_9_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_24_source_9_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_24_source_9_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_24_source_9_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_24_source_9_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_24_source_9_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_24_source_9_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_24_source_9_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_24_source_9_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_24_source_9_pat_stride_buf_3;
  wire _set_flag_407;
  assign _set_flag_407 = conv2d_24_comp_fsm == 3;
  wire [2-1:0] read_rtl_bank_408;
  assign read_rtl_bank_408 = _stream_conv2d_24_source_9_source_ram_raddr;
  reg [2-1:0] _tmp_409;
  localparam _tmp_410 = 1;
  wire [_tmp_410-1:0] _tmp_411;
  assign _tmp_411 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_9_source_ram_renable && (_stream_conv2d_24_source_9_source_sel == 2);
  reg [_tmp_410-1:0] __tmp_411_1;
  localparam _tmp_412 = 1;
  wire [_tmp_412-1:0] _tmp_413;
  assign _tmp_413 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_9_source_ram_renable && (_stream_conv2d_24_source_9_source_sel == 2);
  reg [_tmp_412-1:0] __tmp_413_1;
  localparam _tmp_414 = 1;
  wire [_tmp_414-1:0] _tmp_415;
  assign _tmp_415 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_9_source_ram_renable && (_stream_conv2d_24_source_9_source_sel == 2);
  reg [_tmp_414-1:0] __tmp_415_1;
  localparam _tmp_416 = 1;
  wire [_tmp_416-1:0] _tmp_417;
  assign _tmp_417 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_9_source_ram_renable && (_stream_conv2d_24_source_9_source_sel == 2);
  reg [_tmp_416-1:0] __tmp_417_1;
  wire signed [8-1:0] read_rtl_rdata_418;
  wire read_rtl_rvalid_419;
  assign read_rtl_rdata_418 = (_tmp_409 == 0)? ram_w8_l2048_id0_0_0_rdata : 
                              (_tmp_409 == 1)? ram_w8_l2048_id0_1_0_rdata : 
                              (_tmp_409 == 2)? ram_w8_l2048_id0_2_0_rdata : 
                              (_tmp_409 == 3)? ram_w8_l2048_id0_3_0_rdata : 0;
  assign read_rtl_rvalid_419 = __tmp_411_1;
  assign _stream_conv2d_24_source_9_source_ram_rdata = (_stream_conv2d_24_source_9_source_sel == 2)? read_rtl_rdata_418 : 'hx;
  reg [8-1:0] __variable_wdata_327;
  assign stream_conv2d_24_source_9_data = __variable_wdata_327;
  reg [32-1:0] _stream_conv2d_24_source_9_source_pat_fsm_1;
  localparam _stream_conv2d_24_source_9_source_pat_fsm_1_init = 0;
  wire [32-1:0] _stream_conv2d_24_source_9_source_pat_all_offset;
  assign _stream_conv2d_24_source_9_source_pat_all_offset = _stream_conv2d_24_source_9_source_offset_buf + _source_stream_conv2d_24_source_9_pat_cur_offset_0 + _source_stream_conv2d_24_source_9_pat_cur_offset_1 + _source_stream_conv2d_24_source_9_pat_cur_offset_2 + _source_stream_conv2d_24_source_9_pat_cur_offset_3;
  wire _set_flag_420;
  assign _set_flag_420 = conv2d_24_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_333;
  assign stream_conv2d_24_parameter_10_data = __variable_wdata_333;
  wire _set_flag_421;
  assign _set_flag_421 = conv2d_24_comp_fsm == 3;
  reg [8-1:0] __variable_wdata_334;
  assign stream_conv2d_24_source_11_data = __variable_wdata_334;
  wire _set_flag_422;
  assign _set_flag_422 = conv2d_24_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_340;
  assign stream_conv2d_24_parameter_12_data = __variable_wdata_340;
  wire _set_flag_423;
  assign _set_flag_423 = conv2d_24_comp_fsm == 3;
  reg [8-1:0] __variable_wdata_341;
  assign stream_conv2d_24_source_13_data = __variable_wdata_341;
  wire _set_flag_424;
  assign _set_flag_424 = conv2d_24_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_347;
  assign stream_conv2d_24_parameter_14_data = __variable_wdata_347;
  wire _set_flag_425;
  assign _set_flag_425 = conv2d_24_comp_fsm == 3;
  reg [8-1:0] __variable_wdata_348;
  assign stream_conv2d_24_source_15_data = __variable_wdata_348;
  wire _set_flag_426;
  assign _set_flag_426 = conv2d_24_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_354;
  assign stream_conv2d_24_parameter_16_data = __variable_wdata_354;
  wire _set_flag_427;
  assign _set_flag_427 = conv2d_24_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_355;
  assign stream_conv2d_24_parameter_17_data = __variable_wdata_355;
  wire _set_flag_428;
  assign _set_flag_428 = conv2d_24_comp_fsm == 3;
  reg [5-1:0] __variable_wdata_356;
  assign stream_conv2d_24_parameter_18_data = __variable_wdata_356;
  wire _set_flag_429;
  assign _set_flag_429 = conv2d_24_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_357;
  assign stream_conv2d_24_parameter_19_data = __variable_wdata_357;
  reg [32-1:0] _source_stream_conv2d_24_source_20_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_24_source_20_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_24_source_20_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_24_source_20_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_24_source_20_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_24_source_20_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_24_source_20_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_24_source_20_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_24_source_20_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_24_source_20_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_24_source_20_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_24_source_20_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_24_source_20_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_24_source_20_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_24_source_20_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_24_source_20_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_24_source_20_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_24_source_20_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_24_source_20_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_24_source_20_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_24_source_20_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_24_source_20_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_24_source_20_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_24_source_20_pat_stride_buf_3;
  wire _set_flag_430;
  assign _set_flag_430 = conv2d_24_comp_fsm == 3;
  wire [2-1:0] read_rtl_bank_431;
  assign read_rtl_bank_431 = _stream_conv2d_24_source_20_source_ram_raddr;
  reg [2-1:0] _tmp_432;
  localparam _tmp_433 = 1;
  wire [_tmp_433-1:0] _tmp_434;
  assign _tmp_434 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_20_source_ram_renable && (_stream_conv2d_24_source_20_source_sel == 3);
  reg [_tmp_433-1:0] __tmp_434_1;
  localparam _tmp_435 = 1;
  wire [_tmp_435-1:0] _tmp_436;
  assign _tmp_436 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_20_source_ram_renable && (_stream_conv2d_24_source_20_source_sel == 3);
  reg [_tmp_435-1:0] __tmp_436_1;
  localparam _tmp_437 = 1;
  wire [_tmp_437-1:0] _tmp_438;
  assign _tmp_438 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_20_source_ram_renable && (_stream_conv2d_24_source_20_source_sel == 3);
  reg [_tmp_437-1:0] __tmp_438_1;
  localparam _tmp_439 = 1;
  wire [_tmp_439-1:0] _tmp_440;
  assign _tmp_440 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_20_source_ram_renable && (_stream_conv2d_24_source_20_source_sel == 3);
  reg [_tmp_439-1:0] __tmp_440_1;
  wire signed [8-1:0] read_rtl_rdata_441;
  wire read_rtl_rvalid_442;
  assign read_rtl_rdata_441 = (_tmp_432 == 0)? ram_w8_l16384_id0_0_0_rdata : 
                              (_tmp_432 == 1)? ram_w8_l16384_id0_1_0_rdata : 
                              (_tmp_432 == 2)? ram_w8_l16384_id0_2_0_rdata : 
                              (_tmp_432 == 3)? ram_w8_l16384_id0_3_0_rdata : 0;
  assign read_rtl_rvalid_442 = __tmp_434_1;
  assign _stream_conv2d_24_source_20_source_ram_rdata = (_stream_conv2d_24_source_20_source_sel == 3)? read_rtl_rdata_441 : 'hx;
  reg [8-1:0] __variable_wdata_358;
  assign stream_conv2d_24_source_20_data = __variable_wdata_358;
  reg [32-1:0] _stream_conv2d_24_source_20_source_pat_fsm_2;
  localparam _stream_conv2d_24_source_20_source_pat_fsm_2_init = 0;
  wire [32-1:0] _stream_conv2d_24_source_20_source_pat_all_offset;
  assign _stream_conv2d_24_source_20_source_pat_all_offset = _stream_conv2d_24_source_20_source_offset_buf + _source_stream_conv2d_24_source_20_pat_cur_offset_0 + _source_stream_conv2d_24_source_20_pat_cur_offset_1 + _source_stream_conv2d_24_source_20_pat_cur_offset_2 + _source_stream_conv2d_24_source_20_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_24_source_21_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_24_source_21_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_24_source_21_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_24_source_21_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_24_source_21_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_24_source_21_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_24_source_21_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_24_source_21_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_24_source_21_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_24_source_21_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_24_source_21_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_24_source_21_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_24_source_21_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_24_source_21_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_24_source_21_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_24_source_21_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_24_source_21_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_24_source_21_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_24_source_21_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_24_source_21_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_24_source_21_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_24_source_21_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_24_source_21_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_24_source_21_pat_stride_buf_3;
  wire _set_flag_443;
  assign _set_flag_443 = conv2d_24_comp_fsm == 3;
  wire [2-1:0] read_rtl_bank_444;
  assign read_rtl_bank_444 = _stream_conv2d_24_source_21_source_ram_raddr;
  reg [2-1:0] _tmp_445;
  localparam _tmp_446 = 1;
  wire [_tmp_446-1:0] _tmp_447;
  assign _tmp_447 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_21_source_ram_renable && (_stream_conv2d_24_source_21_source_sel == 4);
  reg [_tmp_446-1:0] __tmp_447_1;
  localparam _tmp_448 = 1;
  wire [_tmp_448-1:0] _tmp_449;
  assign _tmp_449 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_21_source_ram_renable && (_stream_conv2d_24_source_21_source_sel == 4);
  reg [_tmp_448-1:0] __tmp_449_1;
  localparam _tmp_450 = 1;
  wire [_tmp_450-1:0] _tmp_451;
  assign _tmp_451 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_21_source_ram_renable && (_stream_conv2d_24_source_21_source_sel == 4);
  reg [_tmp_450-1:0] __tmp_451_1;
  localparam _tmp_452 = 1;
  wire [_tmp_452-1:0] _tmp_453;
  assign _tmp_453 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_21_source_ram_renable && (_stream_conv2d_24_source_21_source_sel == 4);
  reg [_tmp_452-1:0] __tmp_453_1;
  wire signed [8-1:0] read_rtl_rdata_454;
  wire read_rtl_rvalid_455;
  assign read_rtl_rdata_454 = (_tmp_445 == 0)? ram_w8_l16384_id1_0_0_rdata : 
                              (_tmp_445 == 1)? ram_w8_l16384_id1_1_0_rdata : 
                              (_tmp_445 == 2)? ram_w8_l16384_id1_2_0_rdata : 
                              (_tmp_445 == 3)? ram_w8_l16384_id1_3_0_rdata : 0;
  assign read_rtl_rvalid_455 = __tmp_447_1;
  assign _stream_conv2d_24_source_21_source_ram_rdata = (_stream_conv2d_24_source_21_source_sel == 4)? read_rtl_rdata_454 : 'hx;
  reg [8-1:0] __variable_wdata_359;
  assign stream_conv2d_24_source_21_data = __variable_wdata_359;
  reg [32-1:0] _stream_conv2d_24_source_21_source_pat_fsm_3;
  localparam _stream_conv2d_24_source_21_source_pat_fsm_3_init = 0;
  wire [32-1:0] _stream_conv2d_24_source_21_source_pat_all_offset;
  assign _stream_conv2d_24_source_21_source_pat_all_offset = _stream_conv2d_24_source_21_source_offset_buf + _source_stream_conv2d_24_source_21_pat_cur_offset_0 + _source_stream_conv2d_24_source_21_pat_cur_offset_1 + _source_stream_conv2d_24_source_21_pat_cur_offset_2 + _source_stream_conv2d_24_source_21_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_24_source_22_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_24_source_22_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_24_source_22_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_24_source_22_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_24_source_22_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_24_source_22_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_24_source_22_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_24_source_22_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_24_source_22_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_24_source_22_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_24_source_22_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_24_source_22_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_24_source_22_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_24_source_22_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_24_source_22_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_24_source_22_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_24_source_22_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_24_source_22_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_24_source_22_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_24_source_22_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_24_source_22_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_24_source_22_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_24_source_22_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_24_source_22_pat_stride_buf_3;
  wire _set_flag_456;
  assign _set_flag_456 = conv2d_24_comp_fsm == 3;
  wire [2-1:0] read_rtl_bank_457;
  assign read_rtl_bank_457 = _stream_conv2d_24_source_22_source_ram_raddr;
  reg [2-1:0] _tmp_458;
  assign ram_w8_l16384_id2_0_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_22_source_ram_renable && (_stream_conv2d_24_source_22_source_sel == 5))? _stream_conv2d_24_source_22_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l16384_id2_0_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_22_source_ram_renable && (_stream_conv2d_24_source_22_source_sel == 5))? 1'd1 : 0;
  localparam _tmp_459 = 1;
  wire [_tmp_459-1:0] _tmp_460;
  assign _tmp_460 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_22_source_ram_renable && (_stream_conv2d_24_source_22_source_sel == 5);
  reg [_tmp_459-1:0] __tmp_460_1;
  assign ram_w8_l16384_id2_1_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_22_source_ram_renable && (_stream_conv2d_24_source_22_source_sel == 5))? _stream_conv2d_24_source_22_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l16384_id2_1_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_22_source_ram_renable && (_stream_conv2d_24_source_22_source_sel == 5))? 1'd1 : 0;
  localparam _tmp_461 = 1;
  wire [_tmp_461-1:0] _tmp_462;
  assign _tmp_462 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_22_source_ram_renable && (_stream_conv2d_24_source_22_source_sel == 5);
  reg [_tmp_461-1:0] __tmp_462_1;
  assign ram_w8_l16384_id2_2_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_22_source_ram_renable && (_stream_conv2d_24_source_22_source_sel == 5))? _stream_conv2d_24_source_22_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l16384_id2_2_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_22_source_ram_renable && (_stream_conv2d_24_source_22_source_sel == 5))? 1'd1 : 0;
  localparam _tmp_463 = 1;
  wire [_tmp_463-1:0] _tmp_464;
  assign _tmp_464 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_22_source_ram_renable && (_stream_conv2d_24_source_22_source_sel == 5);
  reg [_tmp_463-1:0] __tmp_464_1;
  assign ram_w8_l16384_id2_3_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_22_source_ram_renable && (_stream_conv2d_24_source_22_source_sel == 5))? _stream_conv2d_24_source_22_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l16384_id2_3_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_22_source_ram_renable && (_stream_conv2d_24_source_22_source_sel == 5))? 1'd1 : 0;
  localparam _tmp_465 = 1;
  wire [_tmp_465-1:0] _tmp_466;
  assign _tmp_466 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_22_source_ram_renable && (_stream_conv2d_24_source_22_source_sel == 5);
  reg [_tmp_465-1:0] __tmp_466_1;
  wire signed [8-1:0] read_rtl_rdata_467;
  wire read_rtl_rvalid_468;
  assign read_rtl_rdata_467 = (_tmp_458 == 0)? ram_w8_l16384_id2_0_0_rdata : 
                              (_tmp_458 == 1)? ram_w8_l16384_id2_1_0_rdata : 
                              (_tmp_458 == 2)? ram_w8_l16384_id2_2_0_rdata : 
                              (_tmp_458 == 3)? ram_w8_l16384_id2_3_0_rdata : 0;
  assign read_rtl_rvalid_468 = __tmp_460_1;
  assign _stream_conv2d_24_source_22_source_ram_rdata = (_stream_conv2d_24_source_22_source_sel == 5)? read_rtl_rdata_467 : 'hx;
  reg [8-1:0] __variable_wdata_360;
  assign stream_conv2d_24_source_22_data = __variable_wdata_360;
  reg [32-1:0] _stream_conv2d_24_source_22_source_pat_fsm_4;
  localparam _stream_conv2d_24_source_22_source_pat_fsm_4_init = 0;
  wire [32-1:0] _stream_conv2d_24_source_22_source_pat_all_offset;
  assign _stream_conv2d_24_source_22_source_pat_all_offset = _stream_conv2d_24_source_22_source_offset_buf + _source_stream_conv2d_24_source_22_pat_cur_offset_0 + _source_stream_conv2d_24_source_22_pat_cur_offset_1 + _source_stream_conv2d_24_source_22_pat_cur_offset_2 + _source_stream_conv2d_24_source_22_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_24_source_23_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_24_source_23_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_24_source_23_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_24_source_23_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_24_source_23_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_24_source_23_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_24_source_23_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_24_source_23_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_24_source_23_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_24_source_23_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_24_source_23_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_24_source_23_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_24_source_23_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_24_source_23_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_24_source_23_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_24_source_23_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_24_source_23_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_24_source_23_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_24_source_23_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_24_source_23_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_24_source_23_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_24_source_23_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_24_source_23_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_24_source_23_pat_stride_buf_3;
  wire _set_flag_469;
  assign _set_flag_469 = conv2d_24_comp_fsm == 3;
  wire [2-1:0] read_rtl_bank_470;
  assign read_rtl_bank_470 = _stream_conv2d_24_source_23_source_ram_raddr;
  reg [2-1:0] _tmp_471;
  assign ram_w8_l16384_id3_0_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_23_source_ram_renable && (_stream_conv2d_24_source_23_source_sel == 6))? _stream_conv2d_24_source_23_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l16384_id3_0_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_23_source_ram_renable && (_stream_conv2d_24_source_23_source_sel == 6))? 1'd1 : 0;
  localparam _tmp_472 = 1;
  wire [_tmp_472-1:0] _tmp_473;
  assign _tmp_473 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_23_source_ram_renable && (_stream_conv2d_24_source_23_source_sel == 6);
  reg [_tmp_472-1:0] __tmp_473_1;
  assign ram_w8_l16384_id3_1_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_23_source_ram_renable && (_stream_conv2d_24_source_23_source_sel == 6))? _stream_conv2d_24_source_23_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l16384_id3_1_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_23_source_ram_renable && (_stream_conv2d_24_source_23_source_sel == 6))? 1'd1 : 0;
  localparam _tmp_474 = 1;
  wire [_tmp_474-1:0] _tmp_475;
  assign _tmp_475 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_23_source_ram_renable && (_stream_conv2d_24_source_23_source_sel == 6);
  reg [_tmp_474-1:0] __tmp_475_1;
  assign ram_w8_l16384_id3_2_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_23_source_ram_renable && (_stream_conv2d_24_source_23_source_sel == 6))? _stream_conv2d_24_source_23_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l16384_id3_2_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_23_source_ram_renable && (_stream_conv2d_24_source_23_source_sel == 6))? 1'd1 : 0;
  localparam _tmp_476 = 1;
  wire [_tmp_476-1:0] _tmp_477;
  assign _tmp_477 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_23_source_ram_renable && (_stream_conv2d_24_source_23_source_sel == 6);
  reg [_tmp_476-1:0] __tmp_477_1;
  assign ram_w8_l16384_id3_3_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_23_source_ram_renable && (_stream_conv2d_24_source_23_source_sel == 6))? _stream_conv2d_24_source_23_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l16384_id3_3_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_23_source_ram_renable && (_stream_conv2d_24_source_23_source_sel == 6))? 1'd1 : 0;
  localparam _tmp_478 = 1;
  wire [_tmp_478-1:0] _tmp_479;
  assign _tmp_479 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_23_source_ram_renable && (_stream_conv2d_24_source_23_source_sel == 6);
  reg [_tmp_478-1:0] __tmp_479_1;
  wire signed [8-1:0] read_rtl_rdata_480;
  wire read_rtl_rvalid_481;
  assign read_rtl_rdata_480 = (_tmp_471 == 0)? ram_w8_l16384_id3_0_0_rdata : 
                              (_tmp_471 == 1)? ram_w8_l16384_id3_1_0_rdata : 
                              (_tmp_471 == 2)? ram_w8_l16384_id3_2_0_rdata : 
                              (_tmp_471 == 3)? ram_w8_l16384_id3_3_0_rdata : 0;
  assign read_rtl_rvalid_481 = __tmp_473_1;
  assign _stream_conv2d_24_source_23_source_ram_rdata = (_stream_conv2d_24_source_23_source_sel == 6)? read_rtl_rdata_480 : 'hx;
  reg [8-1:0] __variable_wdata_361;
  assign stream_conv2d_24_source_23_data = __variable_wdata_361;
  reg [32-1:0] _stream_conv2d_24_source_23_source_pat_fsm_5;
  localparam _stream_conv2d_24_source_23_source_pat_fsm_5_init = 0;
  wire [32-1:0] _stream_conv2d_24_source_23_source_pat_all_offset;
  assign _stream_conv2d_24_source_23_source_pat_all_offset = _stream_conv2d_24_source_23_source_offset_buf + _source_stream_conv2d_24_source_23_pat_cur_offset_0 + _source_stream_conv2d_24_source_23_pat_cur_offset_1 + _source_stream_conv2d_24_source_23_pat_cur_offset_2 + _source_stream_conv2d_24_source_23_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_24_source_24_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_24_source_24_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_24_source_24_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_24_source_24_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_24_source_24_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_24_source_24_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_24_source_24_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_24_source_24_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_24_source_24_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_24_source_24_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_24_source_24_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_24_source_24_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_24_source_24_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_24_source_24_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_24_source_24_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_24_source_24_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_24_source_24_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_24_source_24_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_24_source_24_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_24_source_24_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_24_source_24_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_24_source_24_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_24_source_24_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_24_source_24_pat_stride_buf_3;
  wire _set_flag_482;
  assign _set_flag_482 = conv2d_24_comp_fsm == 3;
  wire [2-1:0] read_rtl_bank_483;
  assign read_rtl_bank_483 = _stream_conv2d_24_source_24_source_ram_raddr;
  reg [2-1:0] _tmp_484;
  assign ram_w8_l16384_id4_0_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_24_source_ram_renable && (_stream_conv2d_24_source_24_source_sel == 7))? _stream_conv2d_24_source_24_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l16384_id4_0_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_24_source_ram_renable && (_stream_conv2d_24_source_24_source_sel == 7))? 1'd1 : 0;
  localparam _tmp_485 = 1;
  wire [_tmp_485-1:0] _tmp_486;
  assign _tmp_486 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_24_source_ram_renable && (_stream_conv2d_24_source_24_source_sel == 7);
  reg [_tmp_485-1:0] __tmp_486_1;
  assign ram_w8_l16384_id4_1_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_24_source_ram_renable && (_stream_conv2d_24_source_24_source_sel == 7))? _stream_conv2d_24_source_24_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l16384_id4_1_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_24_source_ram_renable && (_stream_conv2d_24_source_24_source_sel == 7))? 1'd1 : 0;
  localparam _tmp_487 = 1;
  wire [_tmp_487-1:0] _tmp_488;
  assign _tmp_488 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_24_source_ram_renable && (_stream_conv2d_24_source_24_source_sel == 7);
  reg [_tmp_487-1:0] __tmp_488_1;
  assign ram_w8_l16384_id4_2_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_24_source_ram_renable && (_stream_conv2d_24_source_24_source_sel == 7))? _stream_conv2d_24_source_24_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l16384_id4_2_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_24_source_ram_renable && (_stream_conv2d_24_source_24_source_sel == 7))? 1'd1 : 0;
  localparam _tmp_489 = 1;
  wire [_tmp_489-1:0] _tmp_490;
  assign _tmp_490 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_24_source_ram_renable && (_stream_conv2d_24_source_24_source_sel == 7);
  reg [_tmp_489-1:0] __tmp_490_1;
  assign ram_w8_l16384_id4_3_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_24_source_ram_renable && (_stream_conv2d_24_source_24_source_sel == 7))? _stream_conv2d_24_source_24_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l16384_id4_3_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_24_source_ram_renable && (_stream_conv2d_24_source_24_source_sel == 7))? 1'd1 : 0;
  localparam _tmp_491 = 1;
  wire [_tmp_491-1:0] _tmp_492;
  assign _tmp_492 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_24_source_ram_renable && (_stream_conv2d_24_source_24_source_sel == 7);
  reg [_tmp_491-1:0] __tmp_492_1;
  wire signed [8-1:0] read_rtl_rdata_493;
  wire read_rtl_rvalid_494;
  assign read_rtl_rdata_493 = (_tmp_484 == 0)? ram_w8_l16384_id4_0_0_rdata : 
                              (_tmp_484 == 1)? ram_w8_l16384_id4_1_0_rdata : 
                              (_tmp_484 == 2)? ram_w8_l16384_id4_2_0_rdata : 
                              (_tmp_484 == 3)? ram_w8_l16384_id4_3_0_rdata : 0;
  assign read_rtl_rvalid_494 = __tmp_486_1;
  assign _stream_conv2d_24_source_24_source_ram_rdata = (_stream_conv2d_24_source_24_source_sel == 7)? read_rtl_rdata_493 : 'hx;
  reg [8-1:0] __variable_wdata_362;
  assign stream_conv2d_24_source_24_data = __variable_wdata_362;
  reg [32-1:0] _stream_conv2d_24_source_24_source_pat_fsm_6;
  localparam _stream_conv2d_24_source_24_source_pat_fsm_6_init = 0;
  wire [32-1:0] _stream_conv2d_24_source_24_source_pat_all_offset;
  assign _stream_conv2d_24_source_24_source_pat_all_offset = _stream_conv2d_24_source_24_source_offset_buf + _source_stream_conv2d_24_source_24_pat_cur_offset_0 + _source_stream_conv2d_24_source_24_pat_cur_offset_1 + _source_stream_conv2d_24_source_24_pat_cur_offset_2 + _source_stream_conv2d_24_source_24_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_24_source_25_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_24_source_25_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_24_source_25_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_24_source_25_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_24_source_25_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_24_source_25_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_24_source_25_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_24_source_25_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_24_source_25_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_24_source_25_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_24_source_25_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_24_source_25_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_24_source_25_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_24_source_25_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_24_source_25_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_24_source_25_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_24_source_25_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_24_source_25_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_24_source_25_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_24_source_25_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_24_source_25_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_24_source_25_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_24_source_25_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_24_source_25_pat_stride_buf_3;
  wire _set_flag_495;
  assign _set_flag_495 = conv2d_24_comp_fsm == 3;
  wire [2-1:0] read_rtl_bank_496;
  assign read_rtl_bank_496 = _stream_conv2d_24_source_25_source_ram_raddr;
  reg [2-1:0] _tmp_497;
  assign ram_w8_l16384_id5_0_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_25_source_ram_renable && (_stream_conv2d_24_source_25_source_sel == 8))? _stream_conv2d_24_source_25_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l16384_id5_0_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_25_source_ram_renable && (_stream_conv2d_24_source_25_source_sel == 8))? 1'd1 : 0;
  localparam _tmp_498 = 1;
  wire [_tmp_498-1:0] _tmp_499;
  assign _tmp_499 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_25_source_ram_renable && (_stream_conv2d_24_source_25_source_sel == 8);
  reg [_tmp_498-1:0] __tmp_499_1;
  assign ram_w8_l16384_id5_1_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_25_source_ram_renable && (_stream_conv2d_24_source_25_source_sel == 8))? _stream_conv2d_24_source_25_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l16384_id5_1_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_25_source_ram_renable && (_stream_conv2d_24_source_25_source_sel == 8))? 1'd1 : 0;
  localparam _tmp_500 = 1;
  wire [_tmp_500-1:0] _tmp_501;
  assign _tmp_501 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_25_source_ram_renable && (_stream_conv2d_24_source_25_source_sel == 8);
  reg [_tmp_500-1:0] __tmp_501_1;
  assign ram_w8_l16384_id5_2_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_25_source_ram_renable && (_stream_conv2d_24_source_25_source_sel == 8))? _stream_conv2d_24_source_25_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l16384_id5_2_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_25_source_ram_renable && (_stream_conv2d_24_source_25_source_sel == 8))? 1'd1 : 0;
  localparam _tmp_502 = 1;
  wire [_tmp_502-1:0] _tmp_503;
  assign _tmp_503 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_25_source_ram_renable && (_stream_conv2d_24_source_25_source_sel == 8);
  reg [_tmp_502-1:0] __tmp_503_1;
  assign ram_w8_l16384_id5_3_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_25_source_ram_renable && (_stream_conv2d_24_source_25_source_sel == 8))? _stream_conv2d_24_source_25_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l16384_id5_3_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_25_source_ram_renable && (_stream_conv2d_24_source_25_source_sel == 8))? 1'd1 : 0;
  localparam _tmp_504 = 1;
  wire [_tmp_504-1:0] _tmp_505;
  assign _tmp_505 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_25_source_ram_renable && (_stream_conv2d_24_source_25_source_sel == 8);
  reg [_tmp_504-1:0] __tmp_505_1;
  wire signed [8-1:0] read_rtl_rdata_506;
  wire read_rtl_rvalid_507;
  assign read_rtl_rdata_506 = (_tmp_497 == 0)? ram_w8_l16384_id5_0_0_rdata : 
                              (_tmp_497 == 1)? ram_w8_l16384_id5_1_0_rdata : 
                              (_tmp_497 == 2)? ram_w8_l16384_id5_2_0_rdata : 
                              (_tmp_497 == 3)? ram_w8_l16384_id5_3_0_rdata : 0;
  assign read_rtl_rvalid_507 = __tmp_499_1;
  assign _stream_conv2d_24_source_25_source_ram_rdata = (_stream_conv2d_24_source_25_source_sel == 8)? read_rtl_rdata_506 : 'hx;
  reg [8-1:0] __variable_wdata_363;
  assign stream_conv2d_24_source_25_data = __variable_wdata_363;
  reg [32-1:0] _stream_conv2d_24_source_25_source_pat_fsm_7;
  localparam _stream_conv2d_24_source_25_source_pat_fsm_7_init = 0;
  wire [32-1:0] _stream_conv2d_24_source_25_source_pat_all_offset;
  assign _stream_conv2d_24_source_25_source_pat_all_offset = _stream_conv2d_24_source_25_source_offset_buf + _source_stream_conv2d_24_source_25_pat_cur_offset_0 + _source_stream_conv2d_24_source_25_pat_cur_offset_1 + _source_stream_conv2d_24_source_25_pat_cur_offset_2 + _source_stream_conv2d_24_source_25_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_24_source_26_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_24_source_26_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_24_source_26_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_24_source_26_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_24_source_26_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_24_source_26_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_24_source_26_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_24_source_26_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_24_source_26_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_24_source_26_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_24_source_26_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_24_source_26_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_24_source_26_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_24_source_26_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_24_source_26_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_24_source_26_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_24_source_26_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_24_source_26_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_24_source_26_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_24_source_26_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_24_source_26_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_24_source_26_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_24_source_26_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_24_source_26_pat_stride_buf_3;
  wire _set_flag_508;
  assign _set_flag_508 = conv2d_24_comp_fsm == 3;
  wire [2-1:0] read_rtl_bank_509;
  assign read_rtl_bank_509 = _stream_conv2d_24_source_26_source_ram_raddr;
  reg [2-1:0] _tmp_510;
  assign ram_w8_l16384_id6_0_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_26_source_ram_renable && (_stream_conv2d_24_source_26_source_sel == 9))? _stream_conv2d_24_source_26_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l16384_id6_0_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_26_source_ram_renable && (_stream_conv2d_24_source_26_source_sel == 9))? 1'd1 : 0;
  localparam _tmp_511 = 1;
  wire [_tmp_511-1:0] _tmp_512;
  assign _tmp_512 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_26_source_ram_renable && (_stream_conv2d_24_source_26_source_sel == 9);
  reg [_tmp_511-1:0] __tmp_512_1;
  assign ram_w8_l16384_id6_1_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_26_source_ram_renable && (_stream_conv2d_24_source_26_source_sel == 9))? _stream_conv2d_24_source_26_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l16384_id6_1_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_26_source_ram_renable && (_stream_conv2d_24_source_26_source_sel == 9))? 1'd1 : 0;
  localparam _tmp_513 = 1;
  wire [_tmp_513-1:0] _tmp_514;
  assign _tmp_514 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_26_source_ram_renable && (_stream_conv2d_24_source_26_source_sel == 9);
  reg [_tmp_513-1:0] __tmp_514_1;
  assign ram_w8_l16384_id6_2_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_26_source_ram_renable && (_stream_conv2d_24_source_26_source_sel == 9))? _stream_conv2d_24_source_26_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l16384_id6_2_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_26_source_ram_renable && (_stream_conv2d_24_source_26_source_sel == 9))? 1'd1 : 0;
  localparam _tmp_515 = 1;
  wire [_tmp_515-1:0] _tmp_516;
  assign _tmp_516 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_26_source_ram_renable && (_stream_conv2d_24_source_26_source_sel == 9);
  reg [_tmp_515-1:0] __tmp_516_1;
  assign ram_w8_l16384_id6_3_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_26_source_ram_renable && (_stream_conv2d_24_source_26_source_sel == 9))? _stream_conv2d_24_source_26_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l16384_id6_3_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_26_source_ram_renable && (_stream_conv2d_24_source_26_source_sel == 9))? 1'd1 : 0;
  localparam _tmp_517 = 1;
  wire [_tmp_517-1:0] _tmp_518;
  assign _tmp_518 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_26_source_ram_renable && (_stream_conv2d_24_source_26_source_sel == 9);
  reg [_tmp_517-1:0] __tmp_518_1;
  wire signed [8-1:0] read_rtl_rdata_519;
  wire read_rtl_rvalid_520;
  assign read_rtl_rdata_519 = (_tmp_510 == 0)? ram_w8_l16384_id6_0_0_rdata : 
                              (_tmp_510 == 1)? ram_w8_l16384_id6_1_0_rdata : 
                              (_tmp_510 == 2)? ram_w8_l16384_id6_2_0_rdata : 
                              (_tmp_510 == 3)? ram_w8_l16384_id6_3_0_rdata : 0;
  assign read_rtl_rvalid_520 = __tmp_512_1;
  assign _stream_conv2d_24_source_26_source_ram_rdata = (_stream_conv2d_24_source_26_source_sel == 9)? read_rtl_rdata_519 : 'hx;
  reg [8-1:0] __variable_wdata_364;
  assign stream_conv2d_24_source_26_data = __variable_wdata_364;
  reg [32-1:0] _stream_conv2d_24_source_26_source_pat_fsm_8;
  localparam _stream_conv2d_24_source_26_source_pat_fsm_8_init = 0;
  wire [32-1:0] _stream_conv2d_24_source_26_source_pat_all_offset;
  assign _stream_conv2d_24_source_26_source_pat_all_offset = _stream_conv2d_24_source_26_source_offset_buf + _source_stream_conv2d_24_source_26_pat_cur_offset_0 + _source_stream_conv2d_24_source_26_pat_cur_offset_1 + _source_stream_conv2d_24_source_26_pat_cur_offset_2 + _source_stream_conv2d_24_source_26_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_24_source_27_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_24_source_27_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_24_source_27_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_24_source_27_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_24_source_27_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_24_source_27_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_24_source_27_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_24_source_27_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_24_source_27_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_24_source_27_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_24_source_27_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_24_source_27_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_24_source_27_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_24_source_27_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_24_source_27_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_24_source_27_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_24_source_27_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_24_source_27_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_24_source_27_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_24_source_27_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_24_source_27_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_24_source_27_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_24_source_27_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_24_source_27_pat_stride_buf_3;
  wire _set_flag_521;
  assign _set_flag_521 = conv2d_24_comp_fsm == 3;
  wire [2-1:0] read_rtl_bank_522;
  assign read_rtl_bank_522 = _stream_conv2d_24_source_27_source_ram_raddr;
  reg [2-1:0] _tmp_523;
  assign ram_w8_l16384_id7_0_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_27_source_ram_renable && (_stream_conv2d_24_source_27_source_sel == 10))? _stream_conv2d_24_source_27_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l16384_id7_0_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_27_source_ram_renable && (_stream_conv2d_24_source_27_source_sel == 10))? 1'd1 : 0;
  localparam _tmp_524 = 1;
  wire [_tmp_524-1:0] _tmp_525;
  assign _tmp_525 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_27_source_ram_renable && (_stream_conv2d_24_source_27_source_sel == 10);
  reg [_tmp_524-1:0] __tmp_525_1;
  assign ram_w8_l16384_id7_1_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_27_source_ram_renable && (_stream_conv2d_24_source_27_source_sel == 10))? _stream_conv2d_24_source_27_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l16384_id7_1_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_27_source_ram_renable && (_stream_conv2d_24_source_27_source_sel == 10))? 1'd1 : 0;
  localparam _tmp_526 = 1;
  wire [_tmp_526-1:0] _tmp_527;
  assign _tmp_527 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_27_source_ram_renable && (_stream_conv2d_24_source_27_source_sel == 10);
  reg [_tmp_526-1:0] __tmp_527_1;
  assign ram_w8_l16384_id7_2_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_27_source_ram_renable && (_stream_conv2d_24_source_27_source_sel == 10))? _stream_conv2d_24_source_27_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l16384_id7_2_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_27_source_ram_renable && (_stream_conv2d_24_source_27_source_sel == 10))? 1'd1 : 0;
  localparam _tmp_528 = 1;
  wire [_tmp_528-1:0] _tmp_529;
  assign _tmp_529 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_27_source_ram_renable && (_stream_conv2d_24_source_27_source_sel == 10);
  reg [_tmp_528-1:0] __tmp_529_1;
  assign ram_w8_l16384_id7_3_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_27_source_ram_renable && (_stream_conv2d_24_source_27_source_sel == 10))? _stream_conv2d_24_source_27_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l16384_id7_3_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_27_source_ram_renable && (_stream_conv2d_24_source_27_source_sel == 10))? 1'd1 : 0;
  localparam _tmp_530 = 1;
  wire [_tmp_530-1:0] _tmp_531;
  assign _tmp_531 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_27_source_ram_renable && (_stream_conv2d_24_source_27_source_sel == 10);
  reg [_tmp_530-1:0] __tmp_531_1;
  wire signed [8-1:0] read_rtl_rdata_532;
  wire read_rtl_rvalid_533;
  assign read_rtl_rdata_532 = (_tmp_523 == 0)? ram_w8_l16384_id7_0_0_rdata : 
                              (_tmp_523 == 1)? ram_w8_l16384_id7_1_0_rdata : 
                              (_tmp_523 == 2)? ram_w8_l16384_id7_2_0_rdata : 
                              (_tmp_523 == 3)? ram_w8_l16384_id7_3_0_rdata : 0;
  assign read_rtl_rvalid_533 = __tmp_525_1;
  assign _stream_conv2d_24_source_27_source_ram_rdata = (_stream_conv2d_24_source_27_source_sel == 10)? read_rtl_rdata_532 : 'hx;
  reg [8-1:0] __variable_wdata_365;
  assign stream_conv2d_24_source_27_data = __variable_wdata_365;
  reg [32-1:0] _stream_conv2d_24_source_27_source_pat_fsm_9;
  localparam _stream_conv2d_24_source_27_source_pat_fsm_9_init = 0;
  wire [32-1:0] _stream_conv2d_24_source_27_source_pat_all_offset;
  assign _stream_conv2d_24_source_27_source_pat_all_offset = _stream_conv2d_24_source_27_source_offset_buf + _source_stream_conv2d_24_source_27_pat_cur_offset_0 + _source_stream_conv2d_24_source_27_pat_cur_offset_1 + _source_stream_conv2d_24_source_27_pat_cur_offset_2 + _source_stream_conv2d_24_source_27_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_24_source_28_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_24_source_28_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_24_source_28_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_24_source_28_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_24_source_28_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_24_source_28_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_24_source_28_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_24_source_28_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_24_source_28_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_24_source_28_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_24_source_28_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_24_source_28_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_24_source_28_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_24_source_28_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_24_source_28_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_24_source_28_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_24_source_28_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_24_source_28_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_24_source_28_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_24_source_28_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_24_source_28_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_24_source_28_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_24_source_28_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_24_source_28_pat_stride_buf_3;
  wire _set_flag_534;
  assign _set_flag_534 = conv2d_24_comp_fsm == 3;
  wire [2-1:0] read_rtl_bank_535;
  assign read_rtl_bank_535 = _stream_conv2d_24_source_28_source_ram_raddr;
  reg [2-1:0] _tmp_536;
  assign ram_w8_l16384_id8_0_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_28_source_ram_renable && (_stream_conv2d_24_source_28_source_sel == 11))? _stream_conv2d_24_source_28_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l16384_id8_0_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_28_source_ram_renable && (_stream_conv2d_24_source_28_source_sel == 11))? 1'd1 : 0;
  localparam _tmp_537 = 1;
  wire [_tmp_537-1:0] _tmp_538;
  assign _tmp_538 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_28_source_ram_renable && (_stream_conv2d_24_source_28_source_sel == 11);
  reg [_tmp_537-1:0] __tmp_538_1;
  assign ram_w8_l16384_id8_1_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_28_source_ram_renable && (_stream_conv2d_24_source_28_source_sel == 11))? _stream_conv2d_24_source_28_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l16384_id8_1_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_28_source_ram_renable && (_stream_conv2d_24_source_28_source_sel == 11))? 1'd1 : 0;
  localparam _tmp_539 = 1;
  wire [_tmp_539-1:0] _tmp_540;
  assign _tmp_540 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_28_source_ram_renable && (_stream_conv2d_24_source_28_source_sel == 11);
  reg [_tmp_539-1:0] __tmp_540_1;
  assign ram_w8_l16384_id8_2_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_28_source_ram_renable && (_stream_conv2d_24_source_28_source_sel == 11))? _stream_conv2d_24_source_28_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l16384_id8_2_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_28_source_ram_renable && (_stream_conv2d_24_source_28_source_sel == 11))? 1'd1 : 0;
  localparam _tmp_541 = 1;
  wire [_tmp_541-1:0] _tmp_542;
  assign _tmp_542 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_28_source_ram_renable && (_stream_conv2d_24_source_28_source_sel == 11);
  reg [_tmp_541-1:0] __tmp_542_1;
  assign ram_w8_l16384_id8_3_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_28_source_ram_renable && (_stream_conv2d_24_source_28_source_sel == 11))? _stream_conv2d_24_source_28_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l16384_id8_3_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_28_source_ram_renable && (_stream_conv2d_24_source_28_source_sel == 11))? 1'd1 : 0;
  localparam _tmp_543 = 1;
  wire [_tmp_543-1:0] _tmp_544;
  assign _tmp_544 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_28_source_ram_renable && (_stream_conv2d_24_source_28_source_sel == 11);
  reg [_tmp_543-1:0] __tmp_544_1;
  wire signed [8-1:0] read_rtl_rdata_545;
  wire read_rtl_rvalid_546;
  assign read_rtl_rdata_545 = (_tmp_536 == 0)? ram_w8_l16384_id8_0_0_rdata : 
                              (_tmp_536 == 1)? ram_w8_l16384_id8_1_0_rdata : 
                              (_tmp_536 == 2)? ram_w8_l16384_id8_2_0_rdata : 
                              (_tmp_536 == 3)? ram_w8_l16384_id8_3_0_rdata : 0;
  assign read_rtl_rvalid_546 = __tmp_538_1;
  assign _stream_conv2d_24_source_28_source_ram_rdata = (_stream_conv2d_24_source_28_source_sel == 11)? read_rtl_rdata_545 : 'hx;
  reg [8-1:0] __variable_wdata_366;
  assign stream_conv2d_24_source_28_data = __variable_wdata_366;
  reg [32-1:0] _stream_conv2d_24_source_28_source_pat_fsm_10;
  localparam _stream_conv2d_24_source_28_source_pat_fsm_10_init = 0;
  wire [32-1:0] _stream_conv2d_24_source_28_source_pat_all_offset;
  assign _stream_conv2d_24_source_28_source_pat_all_offset = _stream_conv2d_24_source_28_source_offset_buf + _source_stream_conv2d_24_source_28_pat_cur_offset_0 + _source_stream_conv2d_24_source_28_pat_cur_offset_1 + _source_stream_conv2d_24_source_28_pat_cur_offset_2 + _source_stream_conv2d_24_source_28_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_24_source_29_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_24_source_29_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_24_source_29_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_24_source_29_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_24_source_29_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_24_source_29_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_24_source_29_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_24_source_29_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_24_source_29_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_24_source_29_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_24_source_29_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_24_source_29_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_24_source_29_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_24_source_29_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_24_source_29_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_24_source_29_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_24_source_29_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_24_source_29_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_24_source_29_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_24_source_29_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_24_source_29_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_24_source_29_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_24_source_29_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_24_source_29_pat_stride_buf_3;
  wire _set_flag_547;
  assign _set_flag_547 = conv2d_24_comp_fsm == 3;
  wire [2-1:0] read_rtl_bank_548;
  assign read_rtl_bank_548 = _stream_conv2d_24_source_29_source_ram_raddr;
  reg [2-1:0] _tmp_549;
  assign ram_w8_l4096_id0_0_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_29_source_ram_renable && (_stream_conv2d_24_source_29_source_sel == 12))? _stream_conv2d_24_source_29_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l4096_id0_0_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_29_source_ram_renable && (_stream_conv2d_24_source_29_source_sel == 12))? 1'd1 : 0;
  localparam _tmp_550 = 1;
  wire [_tmp_550-1:0] _tmp_551;
  assign _tmp_551 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_29_source_ram_renable && (_stream_conv2d_24_source_29_source_sel == 12);
  reg [_tmp_550-1:0] __tmp_551_1;
  assign ram_w8_l4096_id0_1_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_29_source_ram_renable && (_stream_conv2d_24_source_29_source_sel == 12))? _stream_conv2d_24_source_29_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l4096_id0_1_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_29_source_ram_renable && (_stream_conv2d_24_source_29_source_sel == 12))? 1'd1 : 0;
  localparam _tmp_552 = 1;
  wire [_tmp_552-1:0] _tmp_553;
  assign _tmp_553 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_29_source_ram_renable && (_stream_conv2d_24_source_29_source_sel == 12);
  reg [_tmp_552-1:0] __tmp_553_1;
  assign ram_w8_l4096_id0_2_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_29_source_ram_renable && (_stream_conv2d_24_source_29_source_sel == 12))? _stream_conv2d_24_source_29_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l4096_id0_2_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_29_source_ram_renable && (_stream_conv2d_24_source_29_source_sel == 12))? 1'd1 : 0;
  localparam _tmp_554 = 1;
  wire [_tmp_554-1:0] _tmp_555;
  assign _tmp_555 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_29_source_ram_renable && (_stream_conv2d_24_source_29_source_sel == 12);
  reg [_tmp_554-1:0] __tmp_555_1;
  assign ram_w8_l4096_id0_3_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_29_source_ram_renable && (_stream_conv2d_24_source_29_source_sel == 12))? _stream_conv2d_24_source_29_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l4096_id0_3_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_29_source_ram_renable && (_stream_conv2d_24_source_29_source_sel == 12))? 1'd1 : 0;
  localparam _tmp_556 = 1;
  wire [_tmp_556-1:0] _tmp_557;
  assign _tmp_557 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_29_source_ram_renable && (_stream_conv2d_24_source_29_source_sel == 12);
  reg [_tmp_556-1:0] __tmp_557_1;
  wire signed [8-1:0] read_rtl_rdata_558;
  wire read_rtl_rvalid_559;
  assign read_rtl_rdata_558 = (_tmp_549 == 0)? ram_w8_l4096_id0_0_0_rdata : 
                              (_tmp_549 == 1)? ram_w8_l4096_id0_1_0_rdata : 
                              (_tmp_549 == 2)? ram_w8_l4096_id0_2_0_rdata : 
                              (_tmp_549 == 3)? ram_w8_l4096_id0_3_0_rdata : 0;
  assign read_rtl_rvalid_559 = __tmp_551_1;
  assign _stream_conv2d_24_source_29_source_ram_rdata = (_stream_conv2d_24_source_29_source_sel == 12)? read_rtl_rdata_558 : 'hx;
  reg [8-1:0] __variable_wdata_592;
  assign stream_conv2d_24_source_29_data = __variable_wdata_592;
  reg [32-1:0] _stream_conv2d_24_source_29_source_pat_fsm_11;
  localparam _stream_conv2d_24_source_29_source_pat_fsm_11_init = 0;
  wire [32-1:0] _stream_conv2d_24_source_29_source_pat_all_offset;
  assign _stream_conv2d_24_source_29_source_pat_all_offset = _stream_conv2d_24_source_29_source_offset_buf + _source_stream_conv2d_24_source_29_pat_cur_offset_0 + _source_stream_conv2d_24_source_29_pat_cur_offset_1 + _source_stream_conv2d_24_source_29_pat_cur_offset_2 + _source_stream_conv2d_24_source_29_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_24_source_30_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_24_source_30_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_24_source_30_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_24_source_30_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_24_source_30_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_24_source_30_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_24_source_30_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_24_source_30_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_24_source_30_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_24_source_30_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_24_source_30_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_24_source_30_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_24_source_30_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_24_source_30_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_24_source_30_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_24_source_30_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_24_source_30_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_24_source_30_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_24_source_30_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_24_source_30_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_24_source_30_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_24_source_30_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_24_source_30_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_24_source_30_pat_stride_buf_3;
  wire _set_flag_560;
  assign _set_flag_560 = conv2d_24_comp_fsm == 3;
  wire [2-1:0] read_rtl_bank_561;
  assign read_rtl_bank_561 = _stream_conv2d_24_source_30_source_ram_raddr;
  reg [2-1:0] _tmp_562;
  assign ram_w8_l4096_id1_0_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_30_source_ram_renable && (_stream_conv2d_24_source_30_source_sel == 13))? _stream_conv2d_24_source_30_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l4096_id1_0_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_30_source_ram_renable && (_stream_conv2d_24_source_30_source_sel == 13))? 1'd1 : 0;
  localparam _tmp_563 = 1;
  wire [_tmp_563-1:0] _tmp_564;
  assign _tmp_564 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_30_source_ram_renable && (_stream_conv2d_24_source_30_source_sel == 13);
  reg [_tmp_563-1:0] __tmp_564_1;
  assign ram_w8_l4096_id1_1_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_30_source_ram_renable && (_stream_conv2d_24_source_30_source_sel == 13))? _stream_conv2d_24_source_30_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l4096_id1_1_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_30_source_ram_renable && (_stream_conv2d_24_source_30_source_sel == 13))? 1'd1 : 0;
  localparam _tmp_565 = 1;
  wire [_tmp_565-1:0] _tmp_566;
  assign _tmp_566 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_30_source_ram_renable && (_stream_conv2d_24_source_30_source_sel == 13);
  reg [_tmp_565-1:0] __tmp_566_1;
  assign ram_w8_l4096_id1_2_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_30_source_ram_renable && (_stream_conv2d_24_source_30_source_sel == 13))? _stream_conv2d_24_source_30_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l4096_id1_2_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_30_source_ram_renable && (_stream_conv2d_24_source_30_source_sel == 13))? 1'd1 : 0;
  localparam _tmp_567 = 1;
  wire [_tmp_567-1:0] _tmp_568;
  assign _tmp_568 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_30_source_ram_renable && (_stream_conv2d_24_source_30_source_sel == 13);
  reg [_tmp_567-1:0] __tmp_568_1;
  assign ram_w8_l4096_id1_3_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_30_source_ram_renable && (_stream_conv2d_24_source_30_source_sel == 13))? _stream_conv2d_24_source_30_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l4096_id1_3_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_30_source_ram_renable && (_stream_conv2d_24_source_30_source_sel == 13))? 1'd1 : 0;
  localparam _tmp_569 = 1;
  wire [_tmp_569-1:0] _tmp_570;
  assign _tmp_570 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_30_source_ram_renable && (_stream_conv2d_24_source_30_source_sel == 13);
  reg [_tmp_569-1:0] __tmp_570_1;
  wire signed [8-1:0] read_rtl_rdata_571;
  wire read_rtl_rvalid_572;
  assign read_rtl_rdata_571 = (_tmp_562 == 0)? ram_w8_l4096_id1_0_0_rdata : 
                              (_tmp_562 == 1)? ram_w8_l4096_id1_1_0_rdata : 
                              (_tmp_562 == 2)? ram_w8_l4096_id1_2_0_rdata : 
                              (_tmp_562 == 3)? ram_w8_l4096_id1_3_0_rdata : 0;
  assign read_rtl_rvalid_572 = __tmp_564_1;
  assign _stream_conv2d_24_source_30_source_ram_rdata = (_stream_conv2d_24_source_30_source_sel == 13)? read_rtl_rdata_571 : 'hx;
  reg [8-1:0] __variable_wdata_593;
  assign stream_conv2d_24_source_30_data = __variable_wdata_593;
  reg [32-1:0] _stream_conv2d_24_source_30_source_pat_fsm_12;
  localparam _stream_conv2d_24_source_30_source_pat_fsm_12_init = 0;
  wire [32-1:0] _stream_conv2d_24_source_30_source_pat_all_offset;
  assign _stream_conv2d_24_source_30_source_pat_all_offset = _stream_conv2d_24_source_30_source_offset_buf + _source_stream_conv2d_24_source_30_pat_cur_offset_0 + _source_stream_conv2d_24_source_30_pat_cur_offset_1 + _source_stream_conv2d_24_source_30_pat_cur_offset_2 + _source_stream_conv2d_24_source_30_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_24_source_31_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_24_source_31_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_24_source_31_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_24_source_31_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_24_source_31_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_24_source_31_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_24_source_31_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_24_source_31_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_24_source_31_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_24_source_31_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_24_source_31_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_24_source_31_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_24_source_31_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_24_source_31_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_24_source_31_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_24_source_31_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_24_source_31_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_24_source_31_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_24_source_31_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_24_source_31_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_24_source_31_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_24_source_31_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_24_source_31_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_24_source_31_pat_stride_buf_3;
  wire _set_flag_573;
  assign _set_flag_573 = conv2d_24_comp_fsm == 3;
  wire [2-1:0] read_rtl_bank_574;
  assign read_rtl_bank_574 = _stream_conv2d_24_source_31_source_ram_raddr;
  reg [2-1:0] _tmp_575;
  assign ram_w8_l4096_id2_0_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_31_source_ram_renable && (_stream_conv2d_24_source_31_source_sel == 14))? _stream_conv2d_24_source_31_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l4096_id2_0_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_31_source_ram_renable && (_stream_conv2d_24_source_31_source_sel == 14))? 1'd1 : 0;
  localparam _tmp_576 = 1;
  wire [_tmp_576-1:0] _tmp_577;
  assign _tmp_577 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_31_source_ram_renable && (_stream_conv2d_24_source_31_source_sel == 14);
  reg [_tmp_576-1:0] __tmp_577_1;
  assign ram_w8_l4096_id2_1_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_31_source_ram_renable && (_stream_conv2d_24_source_31_source_sel == 14))? _stream_conv2d_24_source_31_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l4096_id2_1_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_31_source_ram_renable && (_stream_conv2d_24_source_31_source_sel == 14))? 1'd1 : 0;
  localparam _tmp_578 = 1;
  wire [_tmp_578-1:0] _tmp_579;
  assign _tmp_579 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_31_source_ram_renable && (_stream_conv2d_24_source_31_source_sel == 14);
  reg [_tmp_578-1:0] __tmp_579_1;
  assign ram_w8_l4096_id2_2_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_31_source_ram_renable && (_stream_conv2d_24_source_31_source_sel == 14))? _stream_conv2d_24_source_31_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l4096_id2_2_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_31_source_ram_renable && (_stream_conv2d_24_source_31_source_sel == 14))? 1'd1 : 0;
  localparam _tmp_580 = 1;
  wire [_tmp_580-1:0] _tmp_581;
  assign _tmp_581 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_31_source_ram_renable && (_stream_conv2d_24_source_31_source_sel == 14);
  reg [_tmp_580-1:0] __tmp_581_1;
  assign ram_w8_l4096_id2_3_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_31_source_ram_renable && (_stream_conv2d_24_source_31_source_sel == 14))? _stream_conv2d_24_source_31_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l4096_id2_3_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_31_source_ram_renable && (_stream_conv2d_24_source_31_source_sel == 14))? 1'd1 : 0;
  localparam _tmp_582 = 1;
  wire [_tmp_582-1:0] _tmp_583;
  assign _tmp_583 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_31_source_ram_renable && (_stream_conv2d_24_source_31_source_sel == 14);
  reg [_tmp_582-1:0] __tmp_583_1;
  wire signed [8-1:0] read_rtl_rdata_584;
  wire read_rtl_rvalid_585;
  assign read_rtl_rdata_584 = (_tmp_575 == 0)? ram_w8_l4096_id2_0_0_rdata : 
                              (_tmp_575 == 1)? ram_w8_l4096_id2_1_0_rdata : 
                              (_tmp_575 == 2)? ram_w8_l4096_id2_2_0_rdata : 
                              (_tmp_575 == 3)? ram_w8_l4096_id2_3_0_rdata : 0;
  assign read_rtl_rvalid_585 = __tmp_577_1;
  assign _stream_conv2d_24_source_31_source_ram_rdata = (_stream_conv2d_24_source_31_source_sel == 14)? read_rtl_rdata_584 : 'hx;
  reg [8-1:0] __variable_wdata_594;
  assign stream_conv2d_24_source_31_data = __variable_wdata_594;
  reg [32-1:0] _stream_conv2d_24_source_31_source_pat_fsm_13;
  localparam _stream_conv2d_24_source_31_source_pat_fsm_13_init = 0;
  wire [32-1:0] _stream_conv2d_24_source_31_source_pat_all_offset;
  assign _stream_conv2d_24_source_31_source_pat_all_offset = _stream_conv2d_24_source_31_source_offset_buf + _source_stream_conv2d_24_source_31_pat_cur_offset_0 + _source_stream_conv2d_24_source_31_pat_cur_offset_1 + _source_stream_conv2d_24_source_31_pat_cur_offset_2 + _source_stream_conv2d_24_source_31_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_24_source_32_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_24_source_32_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_24_source_32_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_24_source_32_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_24_source_32_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_24_source_32_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_24_source_32_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_24_source_32_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_24_source_32_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_24_source_32_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_24_source_32_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_24_source_32_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_24_source_32_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_24_source_32_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_24_source_32_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_24_source_32_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_24_source_32_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_24_source_32_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_24_source_32_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_24_source_32_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_24_source_32_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_24_source_32_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_24_source_32_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_24_source_32_pat_stride_buf_3;
  wire _set_flag_586;
  assign _set_flag_586 = conv2d_24_comp_fsm == 3;
  wire [2-1:0] read_rtl_bank_587;
  assign read_rtl_bank_587 = _stream_conv2d_24_source_32_source_ram_raddr;
  reg [2-1:0] _tmp_588;
  assign ram_w8_l4096_id3_0_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_32_source_ram_renable && (_stream_conv2d_24_source_32_source_sel == 15))? _stream_conv2d_24_source_32_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l4096_id3_0_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_32_source_ram_renable && (_stream_conv2d_24_source_32_source_sel == 15))? 1'd1 : 0;
  localparam _tmp_589 = 1;
  wire [_tmp_589-1:0] _tmp_590;
  assign _tmp_590 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_32_source_ram_renable && (_stream_conv2d_24_source_32_source_sel == 15);
  reg [_tmp_589-1:0] __tmp_590_1;
  assign ram_w8_l4096_id3_1_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_32_source_ram_renable && (_stream_conv2d_24_source_32_source_sel == 15))? _stream_conv2d_24_source_32_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l4096_id3_1_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_32_source_ram_renable && (_stream_conv2d_24_source_32_source_sel == 15))? 1'd1 : 0;
  localparam _tmp_591 = 1;
  wire [_tmp_591-1:0] _tmp_592;
  assign _tmp_592 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_32_source_ram_renable && (_stream_conv2d_24_source_32_source_sel == 15);
  reg [_tmp_591-1:0] __tmp_592_1;
  assign ram_w8_l4096_id3_2_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_32_source_ram_renable && (_stream_conv2d_24_source_32_source_sel == 15))? _stream_conv2d_24_source_32_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l4096_id3_2_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_32_source_ram_renable && (_stream_conv2d_24_source_32_source_sel == 15))? 1'd1 : 0;
  localparam _tmp_593 = 1;
  wire [_tmp_593-1:0] _tmp_594;
  assign _tmp_594 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_32_source_ram_renable && (_stream_conv2d_24_source_32_source_sel == 15);
  reg [_tmp_593-1:0] __tmp_594_1;
  assign ram_w8_l4096_id3_3_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_32_source_ram_renable && (_stream_conv2d_24_source_32_source_sel == 15))? _stream_conv2d_24_source_32_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l4096_id3_3_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_32_source_ram_renable && (_stream_conv2d_24_source_32_source_sel == 15))? 1'd1 : 0;
  localparam _tmp_595 = 1;
  wire [_tmp_595-1:0] _tmp_596;
  assign _tmp_596 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_32_source_ram_renable && (_stream_conv2d_24_source_32_source_sel == 15);
  reg [_tmp_595-1:0] __tmp_596_1;
  wire signed [8-1:0] read_rtl_rdata_597;
  wire read_rtl_rvalid_598;
  assign read_rtl_rdata_597 = (_tmp_588 == 0)? ram_w8_l4096_id3_0_0_rdata : 
                              (_tmp_588 == 1)? ram_w8_l4096_id3_1_0_rdata : 
                              (_tmp_588 == 2)? ram_w8_l4096_id3_2_0_rdata : 
                              (_tmp_588 == 3)? ram_w8_l4096_id3_3_0_rdata : 0;
  assign read_rtl_rvalid_598 = __tmp_590_1;
  assign _stream_conv2d_24_source_32_source_ram_rdata = (_stream_conv2d_24_source_32_source_sel == 15)? read_rtl_rdata_597 : 'hx;
  reg [8-1:0] __variable_wdata_595;
  assign stream_conv2d_24_source_32_data = __variable_wdata_595;
  reg [32-1:0] _stream_conv2d_24_source_32_source_pat_fsm_14;
  localparam _stream_conv2d_24_source_32_source_pat_fsm_14_init = 0;
  wire [32-1:0] _stream_conv2d_24_source_32_source_pat_all_offset;
  assign _stream_conv2d_24_source_32_source_pat_all_offset = _stream_conv2d_24_source_32_source_offset_buf + _source_stream_conv2d_24_source_32_pat_cur_offset_0 + _source_stream_conv2d_24_source_32_pat_cur_offset_1 + _source_stream_conv2d_24_source_32_pat_cur_offset_2 + _source_stream_conv2d_24_source_32_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_24_source_33_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_24_source_33_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_24_source_33_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_24_source_33_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_24_source_33_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_24_source_33_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_24_source_33_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_24_source_33_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_24_source_33_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_24_source_33_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_24_source_33_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_24_source_33_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_24_source_33_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_24_source_33_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_24_source_33_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_24_source_33_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_24_source_33_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_24_source_33_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_24_source_33_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_24_source_33_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_24_source_33_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_24_source_33_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_24_source_33_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_24_source_33_pat_stride_buf_3;
  wire _set_flag_599;
  assign _set_flag_599 = conv2d_24_comp_fsm == 3;
  wire [2-1:0] read_rtl_bank_600;
  assign read_rtl_bank_600 = _stream_conv2d_24_source_33_source_ram_raddr;
  reg [2-1:0] _tmp_601;
  assign ram_w8_l4096_id4_0_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_33_source_ram_renable && (_stream_conv2d_24_source_33_source_sel == 16))? _stream_conv2d_24_source_33_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l4096_id4_0_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_33_source_ram_renable && (_stream_conv2d_24_source_33_source_sel == 16))? 1'd1 : 0;
  localparam _tmp_602 = 1;
  wire [_tmp_602-1:0] _tmp_603;
  assign _tmp_603 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_33_source_ram_renable && (_stream_conv2d_24_source_33_source_sel == 16);
  reg [_tmp_602-1:0] __tmp_603_1;
  assign ram_w8_l4096_id4_1_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_33_source_ram_renable && (_stream_conv2d_24_source_33_source_sel == 16))? _stream_conv2d_24_source_33_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l4096_id4_1_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_33_source_ram_renable && (_stream_conv2d_24_source_33_source_sel == 16))? 1'd1 : 0;
  localparam _tmp_604 = 1;
  wire [_tmp_604-1:0] _tmp_605;
  assign _tmp_605 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_33_source_ram_renable && (_stream_conv2d_24_source_33_source_sel == 16);
  reg [_tmp_604-1:0] __tmp_605_1;
  assign ram_w8_l4096_id4_2_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_33_source_ram_renable && (_stream_conv2d_24_source_33_source_sel == 16))? _stream_conv2d_24_source_33_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l4096_id4_2_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_33_source_ram_renable && (_stream_conv2d_24_source_33_source_sel == 16))? 1'd1 : 0;
  localparam _tmp_606 = 1;
  wire [_tmp_606-1:0] _tmp_607;
  assign _tmp_607 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_33_source_ram_renable && (_stream_conv2d_24_source_33_source_sel == 16);
  reg [_tmp_606-1:0] __tmp_607_1;
  assign ram_w8_l4096_id4_3_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_33_source_ram_renable && (_stream_conv2d_24_source_33_source_sel == 16))? _stream_conv2d_24_source_33_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l4096_id4_3_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_33_source_ram_renable && (_stream_conv2d_24_source_33_source_sel == 16))? 1'd1 : 0;
  localparam _tmp_608 = 1;
  wire [_tmp_608-1:0] _tmp_609;
  assign _tmp_609 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_33_source_ram_renable && (_stream_conv2d_24_source_33_source_sel == 16);
  reg [_tmp_608-1:0] __tmp_609_1;
  wire signed [8-1:0] read_rtl_rdata_610;
  wire read_rtl_rvalid_611;
  assign read_rtl_rdata_610 = (_tmp_601 == 0)? ram_w8_l4096_id4_0_0_rdata : 
                              (_tmp_601 == 1)? ram_w8_l4096_id4_1_0_rdata : 
                              (_tmp_601 == 2)? ram_w8_l4096_id4_2_0_rdata : 
                              (_tmp_601 == 3)? ram_w8_l4096_id4_3_0_rdata : 0;
  assign read_rtl_rvalid_611 = __tmp_603_1;
  assign _stream_conv2d_24_source_33_source_ram_rdata = (_stream_conv2d_24_source_33_source_sel == 16)? read_rtl_rdata_610 : 'hx;
  reg [8-1:0] __variable_wdata_596;
  assign stream_conv2d_24_source_33_data = __variable_wdata_596;
  reg [32-1:0] _stream_conv2d_24_source_33_source_pat_fsm_15;
  localparam _stream_conv2d_24_source_33_source_pat_fsm_15_init = 0;
  wire [32-1:0] _stream_conv2d_24_source_33_source_pat_all_offset;
  assign _stream_conv2d_24_source_33_source_pat_all_offset = _stream_conv2d_24_source_33_source_offset_buf + _source_stream_conv2d_24_source_33_pat_cur_offset_0 + _source_stream_conv2d_24_source_33_pat_cur_offset_1 + _source_stream_conv2d_24_source_33_pat_cur_offset_2 + _source_stream_conv2d_24_source_33_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_24_source_34_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_24_source_34_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_24_source_34_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_24_source_34_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_24_source_34_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_24_source_34_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_24_source_34_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_24_source_34_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_24_source_34_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_24_source_34_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_24_source_34_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_24_source_34_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_24_source_34_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_24_source_34_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_24_source_34_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_24_source_34_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_24_source_34_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_24_source_34_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_24_source_34_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_24_source_34_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_24_source_34_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_24_source_34_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_24_source_34_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_24_source_34_pat_stride_buf_3;
  wire _set_flag_612;
  assign _set_flag_612 = conv2d_24_comp_fsm == 3;
  wire [2-1:0] read_rtl_bank_613;
  assign read_rtl_bank_613 = _stream_conv2d_24_source_34_source_ram_raddr;
  reg [2-1:0] _tmp_614;
  assign ram_w8_l4096_id5_0_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_34_source_ram_renable && (_stream_conv2d_24_source_34_source_sel == 17))? _stream_conv2d_24_source_34_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l4096_id5_0_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_34_source_ram_renable && (_stream_conv2d_24_source_34_source_sel == 17))? 1'd1 : 0;
  localparam _tmp_615 = 1;
  wire [_tmp_615-1:0] _tmp_616;
  assign _tmp_616 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_34_source_ram_renable && (_stream_conv2d_24_source_34_source_sel == 17);
  reg [_tmp_615-1:0] __tmp_616_1;
  assign ram_w8_l4096_id5_1_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_34_source_ram_renable && (_stream_conv2d_24_source_34_source_sel == 17))? _stream_conv2d_24_source_34_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l4096_id5_1_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_34_source_ram_renable && (_stream_conv2d_24_source_34_source_sel == 17))? 1'd1 : 0;
  localparam _tmp_617 = 1;
  wire [_tmp_617-1:0] _tmp_618;
  assign _tmp_618 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_34_source_ram_renable && (_stream_conv2d_24_source_34_source_sel == 17);
  reg [_tmp_617-1:0] __tmp_618_1;
  assign ram_w8_l4096_id5_2_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_34_source_ram_renable && (_stream_conv2d_24_source_34_source_sel == 17))? _stream_conv2d_24_source_34_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l4096_id5_2_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_34_source_ram_renable && (_stream_conv2d_24_source_34_source_sel == 17))? 1'd1 : 0;
  localparam _tmp_619 = 1;
  wire [_tmp_619-1:0] _tmp_620;
  assign _tmp_620 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_34_source_ram_renable && (_stream_conv2d_24_source_34_source_sel == 17);
  reg [_tmp_619-1:0] __tmp_620_1;
  assign ram_w8_l4096_id5_3_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_34_source_ram_renable && (_stream_conv2d_24_source_34_source_sel == 17))? _stream_conv2d_24_source_34_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l4096_id5_3_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_34_source_ram_renable && (_stream_conv2d_24_source_34_source_sel == 17))? 1'd1 : 0;
  localparam _tmp_621 = 1;
  wire [_tmp_621-1:0] _tmp_622;
  assign _tmp_622 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_34_source_ram_renable && (_stream_conv2d_24_source_34_source_sel == 17);
  reg [_tmp_621-1:0] __tmp_622_1;
  wire signed [8-1:0] read_rtl_rdata_623;
  wire read_rtl_rvalid_624;
  assign read_rtl_rdata_623 = (_tmp_614 == 0)? ram_w8_l4096_id5_0_0_rdata : 
                              (_tmp_614 == 1)? ram_w8_l4096_id5_1_0_rdata : 
                              (_tmp_614 == 2)? ram_w8_l4096_id5_2_0_rdata : 
                              (_tmp_614 == 3)? ram_w8_l4096_id5_3_0_rdata : 0;
  assign read_rtl_rvalid_624 = __tmp_616_1;
  assign _stream_conv2d_24_source_34_source_ram_rdata = (_stream_conv2d_24_source_34_source_sel == 17)? read_rtl_rdata_623 : 'hx;
  reg [8-1:0] __variable_wdata_597;
  assign stream_conv2d_24_source_34_data = __variable_wdata_597;
  reg [32-1:0] _stream_conv2d_24_source_34_source_pat_fsm_16;
  localparam _stream_conv2d_24_source_34_source_pat_fsm_16_init = 0;
  wire [32-1:0] _stream_conv2d_24_source_34_source_pat_all_offset;
  assign _stream_conv2d_24_source_34_source_pat_all_offset = _stream_conv2d_24_source_34_source_offset_buf + _source_stream_conv2d_24_source_34_pat_cur_offset_0 + _source_stream_conv2d_24_source_34_pat_cur_offset_1 + _source_stream_conv2d_24_source_34_pat_cur_offset_2 + _source_stream_conv2d_24_source_34_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_24_source_35_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_24_source_35_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_24_source_35_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_24_source_35_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_24_source_35_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_24_source_35_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_24_source_35_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_24_source_35_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_24_source_35_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_24_source_35_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_24_source_35_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_24_source_35_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_24_source_35_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_24_source_35_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_24_source_35_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_24_source_35_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_24_source_35_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_24_source_35_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_24_source_35_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_24_source_35_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_24_source_35_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_24_source_35_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_24_source_35_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_24_source_35_pat_stride_buf_3;
  wire _set_flag_625;
  assign _set_flag_625 = conv2d_24_comp_fsm == 3;
  wire [2-1:0] read_rtl_bank_626;
  assign read_rtl_bank_626 = _stream_conv2d_24_source_35_source_ram_raddr;
  reg [2-1:0] _tmp_627;
  assign ram_w8_l4096_id6_0_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_35_source_ram_renable && (_stream_conv2d_24_source_35_source_sel == 18))? _stream_conv2d_24_source_35_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l4096_id6_0_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_35_source_ram_renable && (_stream_conv2d_24_source_35_source_sel == 18))? 1'd1 : 0;
  localparam _tmp_628 = 1;
  wire [_tmp_628-1:0] _tmp_629;
  assign _tmp_629 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_35_source_ram_renable && (_stream_conv2d_24_source_35_source_sel == 18);
  reg [_tmp_628-1:0] __tmp_629_1;
  assign ram_w8_l4096_id6_1_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_35_source_ram_renable && (_stream_conv2d_24_source_35_source_sel == 18))? _stream_conv2d_24_source_35_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l4096_id6_1_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_35_source_ram_renable && (_stream_conv2d_24_source_35_source_sel == 18))? 1'd1 : 0;
  localparam _tmp_630 = 1;
  wire [_tmp_630-1:0] _tmp_631;
  assign _tmp_631 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_35_source_ram_renable && (_stream_conv2d_24_source_35_source_sel == 18);
  reg [_tmp_630-1:0] __tmp_631_1;
  assign ram_w8_l4096_id6_2_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_35_source_ram_renable && (_stream_conv2d_24_source_35_source_sel == 18))? _stream_conv2d_24_source_35_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l4096_id6_2_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_35_source_ram_renable && (_stream_conv2d_24_source_35_source_sel == 18))? 1'd1 : 0;
  localparam _tmp_632 = 1;
  wire [_tmp_632-1:0] _tmp_633;
  assign _tmp_633 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_35_source_ram_renable && (_stream_conv2d_24_source_35_source_sel == 18);
  reg [_tmp_632-1:0] __tmp_633_1;
  assign ram_w8_l4096_id6_3_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_35_source_ram_renable && (_stream_conv2d_24_source_35_source_sel == 18))? _stream_conv2d_24_source_35_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l4096_id6_3_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_35_source_ram_renable && (_stream_conv2d_24_source_35_source_sel == 18))? 1'd1 : 0;
  localparam _tmp_634 = 1;
  wire [_tmp_634-1:0] _tmp_635;
  assign _tmp_635 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_35_source_ram_renable && (_stream_conv2d_24_source_35_source_sel == 18);
  reg [_tmp_634-1:0] __tmp_635_1;
  wire signed [8-1:0] read_rtl_rdata_636;
  wire read_rtl_rvalid_637;
  assign read_rtl_rdata_636 = (_tmp_627 == 0)? ram_w8_l4096_id6_0_0_rdata : 
                              (_tmp_627 == 1)? ram_w8_l4096_id6_1_0_rdata : 
                              (_tmp_627 == 2)? ram_w8_l4096_id6_2_0_rdata : 
                              (_tmp_627 == 3)? ram_w8_l4096_id6_3_0_rdata : 0;
  assign read_rtl_rvalid_637 = __tmp_629_1;
  assign _stream_conv2d_24_source_35_source_ram_rdata = (_stream_conv2d_24_source_35_source_sel == 18)? read_rtl_rdata_636 : 'hx;
  reg [8-1:0] __variable_wdata_598;
  assign stream_conv2d_24_source_35_data = __variable_wdata_598;
  reg [32-1:0] _stream_conv2d_24_source_35_source_pat_fsm_17;
  localparam _stream_conv2d_24_source_35_source_pat_fsm_17_init = 0;
  wire [32-1:0] _stream_conv2d_24_source_35_source_pat_all_offset;
  assign _stream_conv2d_24_source_35_source_pat_all_offset = _stream_conv2d_24_source_35_source_offset_buf + _source_stream_conv2d_24_source_35_pat_cur_offset_0 + _source_stream_conv2d_24_source_35_pat_cur_offset_1 + _source_stream_conv2d_24_source_35_pat_cur_offset_2 + _source_stream_conv2d_24_source_35_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_24_source_36_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_24_source_36_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_24_source_36_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_24_source_36_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_24_source_36_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_24_source_36_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_24_source_36_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_24_source_36_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_24_source_36_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_24_source_36_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_24_source_36_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_24_source_36_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_24_source_36_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_24_source_36_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_24_source_36_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_24_source_36_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_24_source_36_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_24_source_36_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_24_source_36_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_24_source_36_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_24_source_36_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_24_source_36_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_24_source_36_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_24_source_36_pat_stride_buf_3;
  wire _set_flag_638;
  assign _set_flag_638 = conv2d_24_comp_fsm == 3;
  wire [2-1:0] read_rtl_bank_639;
  assign read_rtl_bank_639 = _stream_conv2d_24_source_36_source_ram_raddr;
  reg [2-1:0] _tmp_640;
  assign ram_w8_l4096_id7_0_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_36_source_ram_renable && (_stream_conv2d_24_source_36_source_sel == 19))? _stream_conv2d_24_source_36_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l4096_id7_0_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_36_source_ram_renable && (_stream_conv2d_24_source_36_source_sel == 19))? 1'd1 : 0;
  localparam _tmp_641 = 1;
  wire [_tmp_641-1:0] _tmp_642;
  assign _tmp_642 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_36_source_ram_renable && (_stream_conv2d_24_source_36_source_sel == 19);
  reg [_tmp_641-1:0] __tmp_642_1;
  assign ram_w8_l4096_id7_1_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_36_source_ram_renable && (_stream_conv2d_24_source_36_source_sel == 19))? _stream_conv2d_24_source_36_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l4096_id7_1_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_36_source_ram_renable && (_stream_conv2d_24_source_36_source_sel == 19))? 1'd1 : 0;
  localparam _tmp_643 = 1;
  wire [_tmp_643-1:0] _tmp_644;
  assign _tmp_644 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_36_source_ram_renable && (_stream_conv2d_24_source_36_source_sel == 19);
  reg [_tmp_643-1:0] __tmp_644_1;
  assign ram_w8_l4096_id7_2_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_36_source_ram_renable && (_stream_conv2d_24_source_36_source_sel == 19))? _stream_conv2d_24_source_36_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l4096_id7_2_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_36_source_ram_renable && (_stream_conv2d_24_source_36_source_sel == 19))? 1'd1 : 0;
  localparam _tmp_645 = 1;
  wire [_tmp_645-1:0] _tmp_646;
  assign _tmp_646 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_36_source_ram_renable && (_stream_conv2d_24_source_36_source_sel == 19);
  reg [_tmp_645-1:0] __tmp_646_1;
  assign ram_w8_l4096_id7_3_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_36_source_ram_renable && (_stream_conv2d_24_source_36_source_sel == 19))? _stream_conv2d_24_source_36_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l4096_id7_3_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_36_source_ram_renable && (_stream_conv2d_24_source_36_source_sel == 19))? 1'd1 : 0;
  localparam _tmp_647 = 1;
  wire [_tmp_647-1:0] _tmp_648;
  assign _tmp_648 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_36_source_ram_renable && (_stream_conv2d_24_source_36_source_sel == 19);
  reg [_tmp_647-1:0] __tmp_648_1;
  wire signed [8-1:0] read_rtl_rdata_649;
  wire read_rtl_rvalid_650;
  assign read_rtl_rdata_649 = (_tmp_640 == 0)? ram_w8_l4096_id7_0_0_rdata : 
                              (_tmp_640 == 1)? ram_w8_l4096_id7_1_0_rdata : 
                              (_tmp_640 == 2)? ram_w8_l4096_id7_2_0_rdata : 
                              (_tmp_640 == 3)? ram_w8_l4096_id7_3_0_rdata : 0;
  assign read_rtl_rvalid_650 = __tmp_642_1;
  assign _stream_conv2d_24_source_36_source_ram_rdata = (_stream_conv2d_24_source_36_source_sel == 19)? read_rtl_rdata_649 : 'hx;
  reg [8-1:0] __variable_wdata_599;
  assign stream_conv2d_24_source_36_data = __variable_wdata_599;
  reg [32-1:0] _stream_conv2d_24_source_36_source_pat_fsm_18;
  localparam _stream_conv2d_24_source_36_source_pat_fsm_18_init = 0;
  wire [32-1:0] _stream_conv2d_24_source_36_source_pat_all_offset;
  assign _stream_conv2d_24_source_36_source_pat_all_offset = _stream_conv2d_24_source_36_source_offset_buf + _source_stream_conv2d_24_source_36_pat_cur_offset_0 + _source_stream_conv2d_24_source_36_pat_cur_offset_1 + _source_stream_conv2d_24_source_36_pat_cur_offset_2 + _source_stream_conv2d_24_source_36_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_24_source_37_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_24_source_37_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_24_source_37_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_24_source_37_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_24_source_37_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_24_source_37_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_24_source_37_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_24_source_37_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_24_source_37_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_24_source_37_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_24_source_37_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_24_source_37_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_24_source_37_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_24_source_37_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_24_source_37_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_24_source_37_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_24_source_37_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_24_source_37_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_24_source_37_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_24_source_37_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_24_source_37_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_24_source_37_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_24_source_37_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_24_source_37_pat_stride_buf_3;
  wire _set_flag_651;
  assign _set_flag_651 = conv2d_24_comp_fsm == 3;
  wire [2-1:0] read_rtl_bank_652;
  assign read_rtl_bank_652 = _stream_conv2d_24_source_37_source_ram_raddr;
  reg [2-1:0] _tmp_653;
  assign ram_w8_l4096_id8_0_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_37_source_ram_renable && (_stream_conv2d_24_source_37_source_sel == 20))? _stream_conv2d_24_source_37_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l4096_id8_0_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_37_source_ram_renable && (_stream_conv2d_24_source_37_source_sel == 20))? 1'd1 : 0;
  localparam _tmp_654 = 1;
  wire [_tmp_654-1:0] _tmp_655;
  assign _tmp_655 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_37_source_ram_renable && (_stream_conv2d_24_source_37_source_sel == 20);
  reg [_tmp_654-1:0] __tmp_655_1;
  assign ram_w8_l4096_id8_1_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_37_source_ram_renable && (_stream_conv2d_24_source_37_source_sel == 20))? _stream_conv2d_24_source_37_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l4096_id8_1_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_37_source_ram_renable && (_stream_conv2d_24_source_37_source_sel == 20))? 1'd1 : 0;
  localparam _tmp_656 = 1;
  wire [_tmp_656-1:0] _tmp_657;
  assign _tmp_657 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_37_source_ram_renable && (_stream_conv2d_24_source_37_source_sel == 20);
  reg [_tmp_656-1:0] __tmp_657_1;
  assign ram_w8_l4096_id8_2_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_37_source_ram_renable && (_stream_conv2d_24_source_37_source_sel == 20))? _stream_conv2d_24_source_37_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l4096_id8_2_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_37_source_ram_renable && (_stream_conv2d_24_source_37_source_sel == 20))? 1'd1 : 0;
  localparam _tmp_658 = 1;
  wire [_tmp_658-1:0] _tmp_659;
  assign _tmp_659 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_37_source_ram_renable && (_stream_conv2d_24_source_37_source_sel == 20);
  reg [_tmp_658-1:0] __tmp_659_1;
  assign ram_w8_l4096_id8_3_0_addr = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_37_source_ram_renable && (_stream_conv2d_24_source_37_source_sel == 20))? _stream_conv2d_24_source_37_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l4096_id8_3_0_enable = (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_37_source_ram_renable && (_stream_conv2d_24_source_37_source_sel == 20))? 1'd1 : 0;
  localparam _tmp_660 = 1;
  wire [_tmp_660-1:0] _tmp_661;
  assign _tmp_661 = _stream_conv2d_24_stream_oready && _stream_conv2d_24_source_37_source_ram_renable && (_stream_conv2d_24_source_37_source_sel == 20);
  reg [_tmp_660-1:0] __tmp_661_1;
  wire signed [8-1:0] read_rtl_rdata_662;
  wire read_rtl_rvalid_663;
  assign read_rtl_rdata_662 = (_tmp_653 == 0)? ram_w8_l4096_id8_0_0_rdata : 
                              (_tmp_653 == 1)? ram_w8_l4096_id8_1_0_rdata : 
                              (_tmp_653 == 2)? ram_w8_l4096_id8_2_0_rdata : 
                              (_tmp_653 == 3)? ram_w8_l4096_id8_3_0_rdata : 0;
  assign read_rtl_rvalid_663 = __tmp_655_1;
  assign _stream_conv2d_24_source_37_source_ram_rdata = (_stream_conv2d_24_source_37_source_sel == 20)? read_rtl_rdata_662 : 'hx;
  reg [8-1:0] __variable_wdata_600;
  assign stream_conv2d_24_source_37_data = __variable_wdata_600;
  reg [32-1:0] _stream_conv2d_24_source_37_source_pat_fsm_19;
  localparam _stream_conv2d_24_source_37_source_pat_fsm_19_init = 0;
  wire [32-1:0] _stream_conv2d_24_source_37_source_pat_all_offset;
  assign _stream_conv2d_24_source_37_source_pat_all_offset = _stream_conv2d_24_source_37_source_offset_buf + _source_stream_conv2d_24_source_37_pat_cur_offset_0 + _source_stream_conv2d_24_source_37_pat_cur_offset_1 + _source_stream_conv2d_24_source_37_pat_cur_offset_2 + _source_stream_conv2d_24_source_37_pat_cur_offset_3;
  wire _set_flag_664;
  assign _set_flag_664 = conv2d_24_comp_fsm == 3;
  reg _tmp_665;
  reg _tmp_666;
  reg _tmp_667;
  reg _tmp_668;
  reg _tmp_669;
  reg _tmp_670;
  reg _tmp_671;
  reg _tmp_672;
  reg _tmp_673;
  reg _tmp_674;
  reg _tmp_675;
  reg _tmp_676;
  reg _tmp_677;
  reg _tmp_678;
  reg _tmp_679;
  reg _tmp_680;
  reg _tmp_681;
  reg _tmp_682;
  reg _tmp_683;
  reg _tmp_684;
  reg _tmp_685;
  reg _tmp_686;
  reg _tmp_687;
  reg _tmp_688;
  reg _tmp_689;
  reg _tmp_690;
  reg _tmp_691;
  reg _tmp_692;
  reg _tmp_693;
  reg _tmp_694;
  reg _tmp_695;
  reg _tmp_696;
  reg _tmp_697;
  localparam _tmp_698 = 33;
  wire [_tmp_698-1:0] _tmp_699;
  assign _tmp_699 = conv2d_24_stream_out_local + conv2d_24_out_page_comp_offset_buf;
  reg [_tmp_698-1:0] _tmp_700;
  reg [_tmp_698-1:0] _tmp_701;
  reg [_tmp_698-1:0] _tmp_702;
  reg [_tmp_698-1:0] _tmp_703;
  reg [_tmp_698-1:0] _tmp_704;
  reg [_tmp_698-1:0] _tmp_705;
  reg [_tmp_698-1:0] _tmp_706;
  reg [_tmp_698-1:0] _tmp_707;
  reg [_tmp_698-1:0] _tmp_708;
  reg [_tmp_698-1:0] _tmp_709;
  reg [_tmp_698-1:0] _tmp_710;
  reg [_tmp_698-1:0] _tmp_711;
  reg [_tmp_698-1:0] _tmp_712;
  reg [_tmp_698-1:0] _tmp_713;
  reg [_tmp_698-1:0] _tmp_714;
  reg [_tmp_698-1:0] _tmp_715;
  reg [_tmp_698-1:0] _tmp_716;
  reg [_tmp_698-1:0] _tmp_717;
  reg [_tmp_698-1:0] _tmp_718;
  reg [_tmp_698-1:0] _tmp_719;
  reg [_tmp_698-1:0] _tmp_720;
  reg [_tmp_698-1:0] _tmp_721;
  reg [_tmp_698-1:0] _tmp_722;
  reg [_tmp_698-1:0] _tmp_723;
  reg [_tmp_698-1:0] _tmp_724;
  reg [_tmp_698-1:0] _tmp_725;
  reg [_tmp_698-1:0] _tmp_726;
  reg [_tmp_698-1:0] _tmp_727;
  reg [_tmp_698-1:0] _tmp_728;
  reg [_tmp_698-1:0] _tmp_729;
  reg [_tmp_698-1:0] _tmp_730;
  reg [_tmp_698-1:0] _tmp_731;
  reg [_tmp_698-1:0] _tmp_732;
  reg [32-1:0] _tmp_733;
  reg [32-1:0] _tmp_734;
  reg [32-1:0] _tmp_735;
  reg [32-1:0] _tmp_736;
  reg [32-1:0] _tmp_737;
  reg [32-1:0] _tmp_738;
  reg [32-1:0] _tmp_739;
  reg [32-1:0] _tmp_740;
  reg [32-1:0] _tmp_741;
  reg [32-1:0] _tmp_742;
  reg [32-1:0] _tmp_743;
  reg [32-1:0] _tmp_744;
  reg [32-1:0] _tmp_745;
  reg [32-1:0] _tmp_746;
  reg [32-1:0] _tmp_747;
  reg [32-1:0] _tmp_748;
  reg [32-1:0] _tmp_749;
  reg [32-1:0] _tmp_750;
  reg [32-1:0] _tmp_751;
  reg [32-1:0] _tmp_752;
  reg [32-1:0] _tmp_753;
  reg [32-1:0] _tmp_754;
  reg [32-1:0] _tmp_755;
  reg [32-1:0] _tmp_756;
  reg [32-1:0] _tmp_757;
  reg [32-1:0] _tmp_758;
  reg [32-1:0] _tmp_759;
  reg [32-1:0] _tmp_760;
  reg [32-1:0] _tmp_761;
  reg [32-1:0] _tmp_762;
  reg [32-1:0] _tmp_763;
  reg [32-1:0] _tmp_764;
  reg [32-1:0] _tmp_765;
  wire [2-1:0] write_rtl_bank_766;
  assign write_rtl_bank_766 = _stream_conv2d_24_sink_50_sink_waddr;
  reg [32-1:0] _stream_conv2d_24_sink_50_sink_fsm_20;
  localparam _stream_conv2d_24_sink_50_sink_fsm_20_init = 0;
  wire _set_flag_767;
  assign _set_flag_767 = conv2d_24_comp_fsm == 4;
  assign _stream_conv2d_24_run_flag = (_set_flag_767)? 1 : 0;
  reg _tmp_768;
  reg _tmp_769;
  reg _tmp_770;
  assign _mul_5_source_stop = _mul_5_stream_oready && 1'd0;
  reg _tmp_771;
  reg _tmp_772;
  reg _tmp_773;
  reg _tmp_774;
  reg _tmp_775;
  reg _tmp_776;
  reg _tmp_777;
  reg _tmp_778;
  reg _tmp_779;
  reg _tmp_780;
  assign _mul_5_sink_start = _tmp_780;
  reg _tmp_781;
  reg _tmp_782;
  reg _tmp_783;
  reg _tmp_784;
  reg _tmp_785;
  reg _tmp_786;
  reg _tmp_787;
  reg _tmp_788;
  reg _tmp_789;
  reg _tmp_790;
  assign _mul_5_sink_stop = _tmp_790;
  reg _tmp_791;
  reg _tmp_792;
  reg _tmp_793;
  reg _tmp_794;
  reg _tmp_795;
  reg _tmp_796;
  reg _tmp_797;
  reg _tmp_798;
  reg _tmp_799;
  reg _tmp_800;
  assign _mul_5_sink_busy = _tmp_800;
  reg _tmp_801;
  assign _mul_5_busy = _mul_5_source_busy || _mul_5_sink_busy || _mul_5_busy_reg;
  reg _tmp_802;
  reg _tmp_803;
  reg _tmp_804;
  assign _mul_6_source_stop = _mul_6_stream_oready && 1'd0;
  reg _tmp_805;
  reg _tmp_806;
  reg _tmp_807;
  reg _tmp_808;
  reg _tmp_809;
  reg _tmp_810;
  reg _tmp_811;
  reg _tmp_812;
  reg _tmp_813;
  reg _tmp_814;
  assign _mul_6_sink_start = _tmp_814;
  reg _tmp_815;
  reg _tmp_816;
  reg _tmp_817;
  reg _tmp_818;
  reg _tmp_819;
  reg _tmp_820;
  reg _tmp_821;
  reg _tmp_822;
  reg _tmp_823;
  reg _tmp_824;
  assign _mul_6_sink_stop = _tmp_824;
  reg _tmp_825;
  reg _tmp_826;
  reg _tmp_827;
  reg _tmp_828;
  reg _tmp_829;
  reg _tmp_830;
  reg _tmp_831;
  reg _tmp_832;
  reg _tmp_833;
  reg _tmp_834;
  assign _mul_6_sink_busy = _tmp_834;
  reg _tmp_835;
  assign _mul_6_busy = _mul_6_source_busy || _mul_6_sink_busy || _mul_6_busy_reg;
  reg _tmp_836;
  reg _tmp_837;
  reg _tmp_838;
  assign _mul_7_source_stop = _mul_7_stream_oready && 1'd0;
  reg _tmp_839;
  reg _tmp_840;
  reg _tmp_841;
  reg _tmp_842;
  reg _tmp_843;
  reg _tmp_844;
  reg _tmp_845;
  reg _tmp_846;
  reg _tmp_847;
  reg _tmp_848;
  assign _mul_7_sink_start = _tmp_848;
  reg _tmp_849;
  reg _tmp_850;
  reg _tmp_851;
  reg _tmp_852;
  reg _tmp_853;
  reg _tmp_854;
  reg _tmp_855;
  reg _tmp_856;
  reg _tmp_857;
  reg _tmp_858;
  assign _mul_7_sink_stop = _tmp_858;
  reg _tmp_859;
  reg _tmp_860;
  reg _tmp_861;
  reg _tmp_862;
  reg _tmp_863;
  reg _tmp_864;
  reg _tmp_865;
  reg _tmp_866;
  reg _tmp_867;
  reg _tmp_868;
  assign _mul_7_sink_busy = _tmp_868;
  reg _tmp_869;
  assign _mul_7_busy = _mul_7_source_busy || _mul_7_sink_busy || _mul_7_busy_reg;
  reg _tmp_870;
  reg _tmp_871;
  reg _tmp_872;
  assign _mul_8_source_stop = _mul_8_stream_oready && 1'd0;
  reg _tmp_873;
  reg _tmp_874;
  reg _tmp_875;
  reg _tmp_876;
  reg _tmp_877;
  reg _tmp_878;
  reg _tmp_879;
  reg _tmp_880;
  reg _tmp_881;
  reg _tmp_882;
  assign _mul_8_sink_start = _tmp_882;
  reg _tmp_883;
  reg _tmp_884;
  reg _tmp_885;
  reg _tmp_886;
  reg _tmp_887;
  reg _tmp_888;
  reg _tmp_889;
  reg _tmp_890;
  reg _tmp_891;
  reg _tmp_892;
  assign _mul_8_sink_stop = _tmp_892;
  reg _tmp_893;
  reg _tmp_894;
  reg _tmp_895;
  reg _tmp_896;
  reg _tmp_897;
  reg _tmp_898;
  reg _tmp_899;
  reg _tmp_900;
  reg _tmp_901;
  reg _tmp_902;
  assign _mul_8_sink_busy = _tmp_902;
  reg _tmp_903;
  assign _mul_8_busy = _mul_8_source_busy || _mul_8_sink_busy || _mul_8_busy_reg;
  reg _tmp_904;
  reg _tmp_905;
  reg _tmp_906;
  assign _mul_9_source_stop = _mul_9_stream_oready && 1'd0;
  reg _tmp_907;
  reg _tmp_908;
  reg _tmp_909;
  reg _tmp_910;
  reg _tmp_911;
  reg _tmp_912;
  reg _tmp_913;
  reg _tmp_914;
  reg _tmp_915;
  reg _tmp_916;
  assign _mul_9_sink_start = _tmp_916;
  reg _tmp_917;
  reg _tmp_918;
  reg _tmp_919;
  reg _tmp_920;
  reg _tmp_921;
  reg _tmp_922;
  reg _tmp_923;
  reg _tmp_924;
  reg _tmp_925;
  reg _tmp_926;
  assign _mul_9_sink_stop = _tmp_926;
  reg _tmp_927;
  reg _tmp_928;
  reg _tmp_929;
  reg _tmp_930;
  reg _tmp_931;
  reg _tmp_932;
  reg _tmp_933;
  reg _tmp_934;
  reg _tmp_935;
  reg _tmp_936;
  assign _mul_9_sink_busy = _tmp_936;
  reg _tmp_937;
  assign _mul_9_busy = _mul_9_source_busy || _mul_9_sink_busy || _mul_9_busy_reg;
  reg _tmp_938;
  reg _tmp_939;
  reg _tmp_940;
  assign _mul_10_source_stop = _mul_10_stream_oready && 1'd0;
  reg _tmp_941;
  reg _tmp_942;
  reg _tmp_943;
  reg _tmp_944;
  reg _tmp_945;
  reg _tmp_946;
  reg _tmp_947;
  reg _tmp_948;
  reg _tmp_949;
  reg _tmp_950;
  assign _mul_10_sink_start = _tmp_950;
  reg _tmp_951;
  reg _tmp_952;
  reg _tmp_953;
  reg _tmp_954;
  reg _tmp_955;
  reg _tmp_956;
  reg _tmp_957;
  reg _tmp_958;
  reg _tmp_959;
  reg _tmp_960;
  assign _mul_10_sink_stop = _tmp_960;
  reg _tmp_961;
  reg _tmp_962;
  reg _tmp_963;
  reg _tmp_964;
  reg _tmp_965;
  reg _tmp_966;
  reg _tmp_967;
  reg _tmp_968;
  reg _tmp_969;
  reg _tmp_970;
  assign _mul_10_sink_busy = _tmp_970;
  reg _tmp_971;
  assign _mul_10_busy = _mul_10_source_busy || _mul_10_sink_busy || _mul_10_busy_reg;
  reg _tmp_972;
  reg _tmp_973;
  reg _tmp_974;
  assign _mul_11_source_stop = _mul_11_stream_oready && 1'd0;
  reg _tmp_975;
  reg _tmp_976;
  reg _tmp_977;
  reg _tmp_978;
  reg _tmp_979;
  reg _tmp_980;
  reg _tmp_981;
  reg _tmp_982;
  reg _tmp_983;
  reg _tmp_984;
  assign _mul_11_sink_start = _tmp_984;
  reg _tmp_985;
  reg _tmp_986;
  reg _tmp_987;
  reg _tmp_988;
  reg _tmp_989;
  reg _tmp_990;
  reg _tmp_991;
  reg _tmp_992;
  reg _tmp_993;
  reg _tmp_994;
  assign _mul_11_sink_stop = _tmp_994;
  reg _tmp_995;
  reg _tmp_996;
  reg _tmp_997;
  reg _tmp_998;
  reg _tmp_999;
  reg _tmp_1000;
  reg _tmp_1001;
  reg _tmp_1002;
  reg _tmp_1003;
  reg _tmp_1004;
  assign _mul_11_sink_busy = _tmp_1004;
  reg _tmp_1005;
  assign _mul_11_busy = _mul_11_source_busy || _mul_11_sink_busy || _mul_11_busy_reg;
  reg _tmp_1006;
  reg _tmp_1007;
  reg _tmp_1008;
  assign _mul_12_source_stop = _mul_12_stream_oready && 1'd0;
  reg _tmp_1009;
  reg _tmp_1010;
  reg _tmp_1011;
  reg _tmp_1012;
  reg _tmp_1013;
  reg _tmp_1014;
  reg _tmp_1015;
  reg _tmp_1016;
  reg _tmp_1017;
  reg _tmp_1018;
  assign _mul_12_sink_start = _tmp_1018;
  reg _tmp_1019;
  reg _tmp_1020;
  reg _tmp_1021;
  reg _tmp_1022;
  reg _tmp_1023;
  reg _tmp_1024;
  reg _tmp_1025;
  reg _tmp_1026;
  reg _tmp_1027;
  reg _tmp_1028;
  assign _mul_12_sink_stop = _tmp_1028;
  reg _tmp_1029;
  reg _tmp_1030;
  reg _tmp_1031;
  reg _tmp_1032;
  reg _tmp_1033;
  reg _tmp_1034;
  reg _tmp_1035;
  reg _tmp_1036;
  reg _tmp_1037;
  reg _tmp_1038;
  assign _mul_12_sink_busy = _tmp_1038;
  reg _tmp_1039;
  assign _mul_12_busy = _mul_12_source_busy || _mul_12_sink_busy || _mul_12_busy_reg;
  reg _tmp_1040;
  reg _tmp_1041;
  reg _tmp_1042;
  assign _mul_13_source_stop = _mul_13_stream_oready && 1'd0;
  reg _tmp_1043;
  reg _tmp_1044;
  reg _tmp_1045;
  reg _tmp_1046;
  reg _tmp_1047;
  reg _tmp_1048;
  reg _tmp_1049;
  reg _tmp_1050;
  reg _tmp_1051;
  reg _tmp_1052;
  assign _mul_13_sink_start = _tmp_1052;
  reg _tmp_1053;
  reg _tmp_1054;
  reg _tmp_1055;
  reg _tmp_1056;
  reg _tmp_1057;
  reg _tmp_1058;
  reg _tmp_1059;
  reg _tmp_1060;
  reg _tmp_1061;
  reg _tmp_1062;
  assign _mul_13_sink_stop = _tmp_1062;
  reg _tmp_1063;
  reg _tmp_1064;
  reg _tmp_1065;
  reg _tmp_1066;
  reg _tmp_1067;
  reg _tmp_1068;
  reg _tmp_1069;
  reg _tmp_1070;
  reg _tmp_1071;
  reg _tmp_1072;
  assign _mul_13_sink_busy = _tmp_1072;
  reg _tmp_1073;
  assign _mul_13_busy = _mul_13_source_busy || _mul_13_sink_busy || _mul_13_busy_reg;
  reg _tmp_1074;
  reg _tmp_1075;
  reg _tmp_1076;
  assign _add_tree_3_source_stop = _add_tree_3_stream_oready && 1'd0;
  reg _tmp_1077;
  reg _tmp_1078;
  reg _tmp_1079;
  reg _tmp_1080;
  assign _add_tree_3_sink_start = _tmp_1080;
  reg _tmp_1081;
  reg _tmp_1082;
  reg _tmp_1083;
  reg _tmp_1084;
  assign _add_tree_3_sink_stop = _tmp_1084;
  reg _tmp_1085;
  reg _tmp_1086;
  reg _tmp_1087;
  reg _tmp_1088;
  assign _add_tree_3_sink_busy = _tmp_1088;
  reg _tmp_1089;
  assign _add_tree_3_busy = _add_tree_3_source_busy || _add_tree_3_sink_busy || _add_tree_3_busy_reg;
  reg _tmp_1090;
  reg _tmp_1091;
  reg _tmp_1092;
  reg _tmp_1093;
  reg _tmp_1094;
  reg _tmp_1095;
  reg _tmp_1096;
  reg _tmp_1097;
  reg _tmp_1098;
  reg _tmp_1099;
  assign _acc_1_source_stop = _acc_1_stream_oready && 1'd0;
  reg _tmp_1100;
  reg _tmp_1101;
  reg _tmp_1102;
  reg _tmp_1103;
  reg _tmp_1104;
  reg _tmp_1105;
  reg _tmp_1106;
  assign _acc_1_sink_start = _tmp_1106;
  reg _tmp_1107;
  reg _tmp_1108;
  reg _tmp_1109;
  reg _tmp_1110;
  reg _tmp_1111;
  reg _tmp_1112;
  reg _tmp_1113;
  assign _acc_1_sink_stop = _tmp_1113;
  reg _tmp_1114;
  reg _tmp_1115;
  reg _tmp_1116;
  reg _tmp_1117;
  reg _tmp_1118;
  reg _tmp_1119;
  reg _tmp_1120;
  assign _acc_1_sink_busy = _tmp_1120;
  reg _tmp_1121;
  assign _acc_1_busy = _acc_1_source_busy || _acc_1_sink_busy || _acc_1_busy_reg;
  reg _tmp_1122;
  reg _tmp_1123;
  reg _tmp_1124;
  assign _mul_rshift_round_clip_4_source_stop = _mul_rshift_round_clip_4_stream_oready && 1'd0;
  reg _tmp_1125;
  reg _tmp_1126;
  reg _tmp_1127;
  reg _tmp_1128;
  reg _tmp_1129;
  reg _tmp_1130;
  reg _tmp_1131;
  reg _tmp_1132;
  reg _tmp_1133;
  reg _tmp_1134;
  assign _mul_rshift_round_clip_4_sink_start = _tmp_1134;
  reg _tmp_1135;
  reg _tmp_1136;
  reg _tmp_1137;
  reg _tmp_1138;
  reg _tmp_1139;
  reg _tmp_1140;
  reg _tmp_1141;
  reg _tmp_1142;
  reg _tmp_1143;
  reg _tmp_1144;
  assign _mul_rshift_round_clip_4_sink_stop = _tmp_1144;
  reg _tmp_1145;
  reg _tmp_1146;
  reg _tmp_1147;
  reg _tmp_1148;
  reg _tmp_1149;
  reg _tmp_1150;
  reg _tmp_1151;
  reg _tmp_1152;
  reg _tmp_1153;
  reg _tmp_1154;
  assign _mul_rshift_round_clip_4_sink_busy = _tmp_1154;
  reg _tmp_1155;
  assign _mul_rshift_round_clip_4_busy = _mul_rshift_round_clip_4_source_busy || _mul_rshift_round_clip_4_sink_busy || _mul_rshift_round_clip_4_busy_reg;
  reg _tmp_1156;
  reg _tmp_1157;
  reg _tmp_1158;
  reg _tmp_1159;
  reg _tmp_1160;
  reg _tmp_1161;
  reg [1-1:0] __variable_wdata_309;
  assign stream_conv2d_24__reduce_reset_data = __variable_wdata_309;
  reg _tmp_1162;
  reg _tmp_1163;
  reg _tmp_1164;
  reg _tmp_1165;
  assign _stream_conv2d_24_source_stop = _stream_conv2d_24_stream_oready && (_stream_conv2d_24_source_11_idle && _stream_conv2d_24_source_13_idle && _stream_conv2d_24_source_15_idle && _stream_conv2d_24_source_20_idle && _stream_conv2d_24_source_21_idle && _stream_conv2d_24_source_22_idle && _stream_conv2d_24_source_23_idle && _stream_conv2d_24_source_24_idle && _stream_conv2d_24_source_25_idle && _stream_conv2d_24_source_26_idle && _stream_conv2d_24_source_27_idle && _stream_conv2d_24_source_28_idle && _stream_conv2d_24_source_29_idle && _stream_conv2d_24_source_30_idle && _stream_conv2d_24_source_31_idle && _stream_conv2d_24_source_32_idle && _stream_conv2d_24_source_33_idle && _stream_conv2d_24_source_34_idle && _stream_conv2d_24_source_35_idle && _stream_conv2d_24_source_36_idle && _stream_conv2d_24_source_37_idle && _stream_conv2d_24_source_7_idle && _stream_conv2d_24_source_9_idle && (_stream_conv2d_24_fsm == 3));
  localparam _tmp_1166 = 1;
  wire [_tmp_1166-1:0] _tmp_1167;
  assign _tmp_1167 = _stream_conv2d_24_source_11_idle && _stream_conv2d_24_source_13_idle && _stream_conv2d_24_source_15_idle && _stream_conv2d_24_source_20_idle && _stream_conv2d_24_source_21_idle && _stream_conv2d_24_source_22_idle && _stream_conv2d_24_source_23_idle && _stream_conv2d_24_source_24_idle && _stream_conv2d_24_source_25_idle && _stream_conv2d_24_source_26_idle && _stream_conv2d_24_source_27_idle && _stream_conv2d_24_source_28_idle && _stream_conv2d_24_source_29_idle && _stream_conv2d_24_source_30_idle && _stream_conv2d_24_source_31_idle && _stream_conv2d_24_source_32_idle && _stream_conv2d_24_source_33_idle && _stream_conv2d_24_source_34_idle && _stream_conv2d_24_source_35_idle && _stream_conv2d_24_source_36_idle && _stream_conv2d_24_source_37_idle && _stream_conv2d_24_source_7_idle && _stream_conv2d_24_source_9_idle && (_stream_conv2d_24_fsm == 3);
  reg [_tmp_1166-1:0] _tmp_1168;
  localparam _tmp_1169 = 1;
  wire [_tmp_1169-1:0] _tmp_1170;
  assign _tmp_1170 = _stream_conv2d_24_source_11_idle && _stream_conv2d_24_source_13_idle && _stream_conv2d_24_source_15_idle && _stream_conv2d_24_source_20_idle && _stream_conv2d_24_source_21_idle && _stream_conv2d_24_source_22_idle && _stream_conv2d_24_source_23_idle && _stream_conv2d_24_source_24_idle && _stream_conv2d_24_source_25_idle && _stream_conv2d_24_source_26_idle && _stream_conv2d_24_source_27_idle && _stream_conv2d_24_source_28_idle && _stream_conv2d_24_source_29_idle && _stream_conv2d_24_source_30_idle && _stream_conv2d_24_source_31_idle && _stream_conv2d_24_source_32_idle && _stream_conv2d_24_source_33_idle && _stream_conv2d_24_source_34_idle && _stream_conv2d_24_source_35_idle && _stream_conv2d_24_source_36_idle && _stream_conv2d_24_source_37_idle && _stream_conv2d_24_source_7_idle && _stream_conv2d_24_source_9_idle && (_stream_conv2d_24_fsm == 3);
  reg [_tmp_1169-1:0] _tmp_1171;
  reg _tmp_1172;
  reg _tmp_1173;
  reg _tmp_1174;
  reg _tmp_1175;
  reg _tmp_1176;
  reg _tmp_1177;
  reg _tmp_1178;
  reg _tmp_1179;
  reg _tmp_1180;
  reg _tmp_1181;
  reg _tmp_1182;
  reg _tmp_1183;
  reg _tmp_1184;
  reg _tmp_1185;
  reg _tmp_1186;
  reg _tmp_1187;
  reg _tmp_1188;
  reg _tmp_1189;
  reg _tmp_1190;
  reg _tmp_1191;
  reg _tmp_1192;
  reg _tmp_1193;
  reg _tmp_1194;
  reg _tmp_1195;
  reg _tmp_1196;
  reg _tmp_1197;
  reg _tmp_1198;
  reg _tmp_1199;
  reg _tmp_1200;
  reg _tmp_1201;
  reg _tmp_1202;
  reg _tmp_1203;
  reg _tmp_1204;
  assign _stream_conv2d_24_sink_start = _tmp_1204;
  reg _tmp_1205;
  reg _tmp_1206;
  reg _tmp_1207;
  reg _tmp_1208;
  reg _tmp_1209;
  reg _tmp_1210;
  reg _tmp_1211;
  reg _tmp_1212;
  reg _tmp_1213;
  reg _tmp_1214;
  reg _tmp_1215;
  reg _tmp_1216;
  reg _tmp_1217;
  reg _tmp_1218;
  reg _tmp_1219;
  reg _tmp_1220;
  reg _tmp_1221;
  reg _tmp_1222;
  reg _tmp_1223;
  reg _tmp_1224;
  reg _tmp_1225;
  reg _tmp_1226;
  reg _tmp_1227;
  reg _tmp_1228;
  reg _tmp_1229;
  reg _tmp_1230;
  reg _tmp_1231;
  reg _tmp_1232;
  reg _tmp_1233;
  reg _tmp_1234;
  reg _tmp_1235;
  reg _tmp_1236;
  reg _tmp_1237;
  assign _stream_conv2d_24_sink_stop = _tmp_1237;
  reg _tmp_1238;
  reg _tmp_1239;
  reg _tmp_1240;
  reg _tmp_1241;
  reg _tmp_1242;
  reg _tmp_1243;
  reg _tmp_1244;
  reg _tmp_1245;
  reg _tmp_1246;
  reg _tmp_1247;
  reg _tmp_1248;
  reg _tmp_1249;
  reg _tmp_1250;
  reg _tmp_1251;
  reg _tmp_1252;
  reg _tmp_1253;
  reg _tmp_1254;
  reg _tmp_1255;
  reg _tmp_1256;
  reg _tmp_1257;
  reg _tmp_1258;
  reg _tmp_1259;
  reg _tmp_1260;
  reg _tmp_1261;
  reg _tmp_1262;
  reg _tmp_1263;
  reg _tmp_1264;
  reg _tmp_1265;
  reg _tmp_1266;
  reg _tmp_1267;
  reg _tmp_1268;
  reg _tmp_1269;
  reg _tmp_1270;
  assign _stream_conv2d_24_sink_busy = _tmp_1270;
  reg _tmp_1271;
  assign _stream_conv2d_24_busy = _stream_conv2d_24_source_busy || _stream_conv2d_24_sink_busy || _stream_conv2d_24_busy_reg;
  wire conv2d_24_dma_out_mask_0;
  assign conv2d_24_dma_out_mask_0 = conv2d_24_out_row_count + 0 >= cparam_conv2d_24_out_num_row;
  wire [32-1:0] _dma_write_packed_high_local_size_1272;
  assign _dma_write_packed_high_local_size_1272 = conv2d_24_next_out_write_size >> 2;
  wire [2-1:0] _dma_write_packed_low_local_size_1273;
  assign _dma_write_packed_low_local_size_1273 = conv2d_24_next_out_write_size & { 2{ 1'd1 } };
  wire [32-1:0] _dma_write_packed_local_packed_size_1274;
  assign _dma_write_packed_local_packed_size_1274 = (_dma_write_packed_low_local_size_1273 > 0)? _dma_write_packed_high_local_size_1272 + 1 : _dma_write_packed_high_local_size_1272;
  wire [32-1:0] mask_addr_shifted_1275;
  assign mask_addr_shifted_1275 = conv2d_24_objaddr + (conv2d_24_out_base_offset + cparam_conv2d_24_out_offset_values_0) + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_1276;
  assign mask_addr_masked_1276 = mask_addr_shifted_1275 << 2;
  reg [32-1:0] _maxi_write_req_fsm;
  localparam _maxi_write_req_fsm_init = 0;
  reg [33-1:0] _maxi_write_cur_global_size;
  reg _maxi_write_cont;
  wire [8-1:0] pack_write_req_op_sel_1277;
  wire [32-1:0] pack_write_req_local_addr_1278;
  wire [32-1:0] pack_write_req_local_stride_1279;
  wire [33-1:0] pack_write_req_size_1280;
  wire [32-1:0] pack_write_req_local_blocksize_1281;
  assign pack_write_req_op_sel_1277 = _maxi_write_op_sel;
  assign pack_write_req_local_addr_1278 = _maxi_write_local_addr;
  assign pack_write_req_local_stride_1279 = _maxi_write_local_stride;
  assign pack_write_req_size_1280 = _maxi_write_local_size;
  assign pack_write_req_local_blocksize_1281 = _maxi_write_local_blocksize;
  wire [137-1:0] pack_write_req_packed_1282;
  assign pack_write_req_packed_1282 = { pack_write_req_op_sel_1277, pack_write_req_local_addr_1278, pack_write_req_local_stride_1279, pack_write_req_size_1280, pack_write_req_local_blocksize_1281 };
  localparam _tmp_1283 = 1;
  wire [_tmp_1283-1:0] _tmp_1284;
  assign _tmp_1284 = !_maxi_write_req_fifo_almost_full;
  reg [_tmp_1283-1:0] __tmp_1284_1;
  wire [32-1:0] mask_addr_shifted_1285;
  assign mask_addr_shifted_1285 = _maxi_write_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_1286;
  assign mask_addr_masked_1286 = mask_addr_shifted_1285 << 2;
  wire [32-1:0] mask_addr_shifted_1287;
  assign mask_addr_shifted_1287 = _maxi_write_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_1288;
  assign mask_addr_masked_1288 = mask_addr_shifted_1287 << 2;
  wire [32-1:0] mask_addr_shifted_1289;
  assign mask_addr_shifted_1289 = _maxi_write_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_1290;
  assign mask_addr_masked_1290 = mask_addr_shifted_1289 << 2;
  wire [32-1:0] mask_addr_shifted_1291;
  assign mask_addr_shifted_1291 = _maxi_write_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_1292;
  assign mask_addr_masked_1292 = mask_addr_shifted_1291 << 2;
  wire [32-1:0] mask_addr_shifted_1293;
  assign mask_addr_shifted_1293 = _maxi_write_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_1294;
  assign mask_addr_masked_1294 = mask_addr_shifted_1293 << 2;
  wire [32-1:0] mask_addr_shifted_1295;
  assign mask_addr_shifted_1295 = _maxi_write_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_1296;
  assign mask_addr_masked_1296 = mask_addr_shifted_1295 << 2;
  wire [8-1:0] pack_write_req_op_sel_1297;
  wire [32-1:0] pack_write_req_local_addr_1298;
  wire [32-1:0] pack_write_req_local_stride_1299;
  wire [33-1:0] pack_write_req_size_1300;
  wire [32-1:0] pack_write_req_local_blocksize_1301;
  assign pack_write_req_op_sel_1297 = _maxi_write_op_sel;
  assign pack_write_req_local_addr_1298 = _maxi_write_local_addr;
  assign pack_write_req_local_stride_1299 = _maxi_write_local_stride;
  assign pack_write_req_size_1300 = _maxi_write_cur_global_size;
  assign pack_write_req_local_blocksize_1301 = _maxi_write_local_blocksize;
  wire [137-1:0] pack_write_req_packed_1302;
  assign pack_write_req_packed_1302 = { pack_write_req_op_sel_1297, pack_write_req_local_addr_1298, pack_write_req_local_stride_1299, pack_write_req_size_1300, pack_write_req_local_blocksize_1301 };
  assign _maxi_write_req_fifo_wdata = ((_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (maxi_awready || !maxi_awvalid) && (_maxi_outstanding_wcount < 6))? pack_write_req_packed_1302 : 
                                      ((_maxi_write_req_fsm == 0) && _maxi_write_start && !_maxi_write_req_fifo_almost_full)? pack_write_req_packed_1282 : 'hx;
  assign _maxi_write_req_fifo_enq = ((_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (maxi_awready || !maxi_awvalid) && (_maxi_outstanding_wcount < 6))? (_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (maxi_awready || !maxi_awvalid) && (_maxi_outstanding_wcount < 6) && !_maxi_write_req_fifo_almost_full : 
                                    ((_maxi_write_req_fsm == 0) && _maxi_write_start && !_maxi_write_req_fifo_almost_full)? (_maxi_write_req_fsm == 0) && _maxi_write_start && !_maxi_write_req_fifo_almost_full && !_maxi_write_req_fifo_almost_full : 0;
  localparam _tmp_1303 = 1;
  wire [_tmp_1303-1:0] _tmp_1304;
  assign _tmp_1304 = !_maxi_write_req_fifo_almost_full;
  reg [_tmp_1303-1:0] __tmp_1304_1;
  reg _maxi_waddr_cond_0_1;
  reg [32-1:0] _maxi_write_data_fsm;
  localparam _maxi_write_data_fsm_init = 0;
  reg [32-1:0] read_burst_packed_fsm_24;
  localparam read_burst_packed_fsm_24_init = 0;
  reg [11-1:0] read_burst_packed_addr_1305;
  reg [11-1:0] read_burst_packed_stride_1306;
  reg [33-1:0] read_burst_packed_length_1307;
  reg read_burst_packed_rvalid_1308;
  reg read_burst_packed_rlast_1309;
  wire [9-1:0] read_burst_packed_ram_addr_1310;
  assign read_burst_packed_ram_addr_1310 = read_burst_packed_addr_1305 >> 2;
  assign ram_w8_l2048_id1_0_1_addr = ((read_burst_packed_fsm_24 == 1) && (!read_burst_packed_rvalid_1308 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)))? read_burst_packed_ram_addr_1310 : 'hx;
  assign ram_w8_l2048_id1_0_1_enable = ((read_burst_packed_fsm_24 == 1) && (!read_burst_packed_rvalid_1308 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)))? 1'd1 : 0;
  localparam _tmp_1311 = 1;
  wire [_tmp_1311-1:0] _tmp_1312;
  assign _tmp_1312 = (read_burst_packed_fsm_24 == 1) && (!read_burst_packed_rvalid_1308 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0));
  reg [_tmp_1311-1:0] __tmp_1312_1;
  wire [8-1:0] read_burst_packed_ram_rdata_1313;
  assign read_burst_packed_ram_rdata_1313 = ram_w8_l2048_id1_0_1_rdata;
  wire [9-1:0] read_burst_packed_ram_addr_1314;
  assign read_burst_packed_ram_addr_1314 = read_burst_packed_addr_1305 >> 2;
  assign ram_w8_l2048_id1_1_1_addr = ((read_burst_packed_fsm_24 == 1) && (!read_burst_packed_rvalid_1308 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)))? read_burst_packed_ram_addr_1314 : 'hx;
  assign ram_w8_l2048_id1_1_1_enable = ((read_burst_packed_fsm_24 == 1) && (!read_burst_packed_rvalid_1308 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)))? 1'd1 : 0;
  localparam _tmp_1315 = 1;
  wire [_tmp_1315-1:0] _tmp_1316;
  assign _tmp_1316 = (read_burst_packed_fsm_24 == 1) && (!read_burst_packed_rvalid_1308 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0));
  reg [_tmp_1315-1:0] __tmp_1316_1;
  wire [8-1:0] read_burst_packed_ram_rdata_1317;
  assign read_burst_packed_ram_rdata_1317 = ram_w8_l2048_id1_1_1_rdata;
  wire [9-1:0] read_burst_packed_ram_addr_1318;
  assign read_burst_packed_ram_addr_1318 = read_burst_packed_addr_1305 >> 2;
  assign ram_w8_l2048_id1_2_1_addr = ((read_burst_packed_fsm_24 == 1) && (!read_burst_packed_rvalid_1308 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)))? read_burst_packed_ram_addr_1318 : 'hx;
  assign ram_w8_l2048_id1_2_1_enable = ((read_burst_packed_fsm_24 == 1) && (!read_burst_packed_rvalid_1308 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)))? 1'd1 : 0;
  localparam _tmp_1319 = 1;
  wire [_tmp_1319-1:0] _tmp_1320;
  assign _tmp_1320 = (read_burst_packed_fsm_24 == 1) && (!read_burst_packed_rvalid_1308 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0));
  reg [_tmp_1319-1:0] __tmp_1320_1;
  wire [8-1:0] read_burst_packed_ram_rdata_1321;
  assign read_burst_packed_ram_rdata_1321 = ram_w8_l2048_id1_2_1_rdata;
  wire [9-1:0] read_burst_packed_ram_addr_1322;
  assign read_burst_packed_ram_addr_1322 = read_burst_packed_addr_1305 >> 2;
  assign ram_w8_l2048_id1_3_1_addr = ((read_burst_packed_fsm_24 == 1) && (!read_burst_packed_rvalid_1308 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)))? read_burst_packed_ram_addr_1322 : 'hx;
  assign ram_w8_l2048_id1_3_1_enable = ((read_burst_packed_fsm_24 == 1) && (!read_burst_packed_rvalid_1308 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)))? 1'd1 : 0;
  localparam _tmp_1323 = 1;
  wire [_tmp_1323-1:0] _tmp_1324;
  assign _tmp_1324 = (read_burst_packed_fsm_24 == 1) && (!read_burst_packed_rvalid_1308 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0));
  reg [_tmp_1323-1:0] __tmp_1324_1;
  wire [8-1:0] read_burst_packed_ram_rdata_1325;
  assign read_burst_packed_ram_rdata_1325 = ram_w8_l2048_id1_3_1_rdata;
  wire [32-1:0] read_burst_packed_rdata_1326;
  assign read_burst_packed_rdata_1326 = { read_burst_packed_ram_rdata_1325, read_burst_packed_ram_rdata_1321, read_burst_packed_ram_rdata_1317, read_burst_packed_ram_rdata_1313 };
  reg _maxi_wdata_cond_0_1;
  wire conv2d_24_update_filter;
  assign conv2d_24_update_filter = (cparam_conv2d_24_data_stationary == 0) && (conv2d_24_row_count >= cparam_conv2d_24_max_row_count) && (conv2d_24_bat_count >= cparam_conv2d_24_max_bat_count) || (cparam_conv2d_24_data_stationary == 1) && !cparam_conv2d_24_keep_filter;
  wire conv2d_24_update_act;
  assign conv2d_24_update_act = (cparam_conv2d_24_data_stationary == 1) && (conv2d_24_och_count >= cparam_conv2d_24_max_och_count) || (cparam_conv2d_24_data_stationary == 0);
  wire conv2d_24_mux_next_dma_flag_0;
  assign conv2d_24_mux_next_dma_flag_0 = (conv2d_24_row_select == 0)? (conv2d_24_row_count >= cparam_conv2d_24_max_row_count)? 1 : cparam_conv2d_24_dma_flag_conds_0 : 
                                         (conv2d_24_row_select == 1)? (conv2d_24_row_count >= cparam_conv2d_24_max_row_count)? 1 : cparam_conv2d_24_dma_flag_conds_2 : 
                                         (conv2d_24_row_select == 2)? (conv2d_24_row_count >= cparam_conv2d_24_max_row_count)? 1 : cparam_conv2d_24_dma_flag_conds_1 : 1'd0;
  wire conv2d_24_mux_next_dma_flag_1;
  assign conv2d_24_mux_next_dma_flag_1 = (conv2d_24_row_select == 0)? (conv2d_24_row_count >= cparam_conv2d_24_max_row_count)? 1 : cparam_conv2d_24_dma_flag_conds_1 : 
                                         (conv2d_24_row_select == 1)? (conv2d_24_row_count >= cparam_conv2d_24_max_row_count)? 1 : cparam_conv2d_24_dma_flag_conds_0 : 
                                         (conv2d_24_row_select == 2)? (conv2d_24_row_count >= cparam_conv2d_24_max_row_count)? 1 : cparam_conv2d_24_dma_flag_conds_2 : 1'd0;
  wire conv2d_24_mux_next_dma_flag_2;
  assign conv2d_24_mux_next_dma_flag_2 = (conv2d_24_row_select == 0)? (conv2d_24_row_count >= cparam_conv2d_24_max_row_count)? 1 : cparam_conv2d_24_dma_flag_conds_2 : 
                                         (conv2d_24_row_select == 1)? (conv2d_24_row_count >= cparam_conv2d_24_max_row_count)? 1 : cparam_conv2d_24_dma_flag_conds_1 : 
                                         (conv2d_24_row_select == 2)? (conv2d_24_row_count >= cparam_conv2d_24_max_row_count)? 1 : cparam_conv2d_24_dma_flag_conds_0 : 1'd0;
  reg [32-1:0] max_pool_serial_26_objaddr;
  reg [32-1:0] max_pool_serial_26_arg_objaddr_0;
  reg [32-1:0] control_max_pool_serial_26;
  localparam control_max_pool_serial_26_init = 0;
  reg _control_max_pool_serial_26_called;
  wire signed [32-1:0] max_pool_serial_26_act_base_offset;
  reg signed [32-1:0] max_pool_serial_26_act_base_offset_row;
  reg signed [32-1:0] max_pool_serial_26_act_base_offset_bat;
  assign max_pool_serial_26_act_base_offset = max_pool_serial_26_act_base_offset_row + max_pool_serial_26_act_base_offset_bat;
  wire signed [32-1:0] max_pool_serial_26_out_base_offset;
  reg signed [32-1:0] max_pool_serial_26_out_base_offset_row;
  reg signed [32-1:0] max_pool_serial_26_out_base_offset_bat;
  assign max_pool_serial_26_out_base_offset = max_pool_serial_26_out_base_offset_row + max_pool_serial_26_out_base_offset_bat;
  reg [32-1:0] max_pool_serial_26_col_count;
  reg [32-1:0] max_pool_serial_26_row_count;
  reg [32-1:0] max_pool_serial_26_bat_count;
  reg [32-1:0] max_pool_serial_26_prev_row_count;
  reg [32-1:0] max_pool_serial_26_prev_bat_count;
  reg [32-1:0] max_pool_serial_26_stream_act_local;
  reg [32-1:0] max_pool_serial_26_stream_out_local;
  reg max_pool_serial_26_act_page;
  reg [32-1:0] max_pool_serial_26_act_page_comp_offset;
  reg [32-1:0] max_pool_serial_26_act_page_dma_offset;
  reg max_pool_serial_26_out_page;
  reg [32-1:0] max_pool_serial_26_out_page_comp_offset;
  reg [32-1:0] max_pool_serial_26_out_page_dma_offset;
  reg max_pool_serial_26_skip_read_act;
  reg max_pool_serial_26_skip_comp;
  reg max_pool_serial_26_skip_write_out;
  reg [32-1:0] max_pool_serial_26_comp_count;
  reg [32-1:0] max_pool_serial_26_out_count;
  wire max_pool_serial_26_dma_pad_mask_0;
  assign max_pool_serial_26_dma_pad_mask_0 = (max_pool_serial_26_row_count + 0 < cparam_max_pool_serial_26_pad_row_top) || (max_pool_serial_26_row_count + 0 >= cparam_max_pool_serial_26_act_num_row + cparam_max_pool_serial_26_pad_row_top);
  wire max_pool_serial_26_dma_pad_mask_1;
  assign max_pool_serial_26_dma_pad_mask_1 = (max_pool_serial_26_row_count + 1 < cparam_max_pool_serial_26_pad_row_top) || (max_pool_serial_26_row_count + 1 >= cparam_max_pool_serial_26_act_num_row + cparam_max_pool_serial_26_pad_row_top);
  wire [14-1:0] _dma_read_packed_high_local_size_1327;
  assign _dma_read_packed_high_local_size_1327 = cparam_max_pool_serial_26_act_read_size >> 2;
  wire [2-1:0] _dma_read_packed_low_local_size_1328;
  assign _dma_read_packed_low_local_size_1328 = cparam_max_pool_serial_26_act_read_size & { 2{ 1'd1 } };
  wire [14-1:0] _dma_read_packed_local_packed_size_1329;
  assign _dma_read_packed_local_packed_size_1329 = (_dma_read_packed_low_local_size_1328 > 0)? _dma_read_packed_high_local_size_1327 + 1 : _dma_read_packed_high_local_size_1327;
  wire [32-1:0] mask_addr_shifted_1330;
  assign mask_addr_shifted_1330 = max_pool_serial_26_arg_objaddr_0 + (max_pool_serial_26_act_base_offset + cparam_max_pool_serial_26_act_offset_values_0) + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_1331;
  assign mask_addr_masked_1331 = mask_addr_shifted_1330 << 2;
  reg [32-1:0] write_burst_packed_fsm_25;
  localparam write_burst_packed_fsm_25_init = 0;
  reg [18-1:0] write_burst_packed_addr_1332;
  reg [18-1:0] write_burst_packed_stride_1333;
  reg [33-1:0] write_burst_packed_length_1334;
  reg write_burst_packed_done_1335;
  wire [16-1:0] write_burst_packed_ram_addr_1336;
  assign write_burst_packed_ram_addr_1336 = write_burst_packed_addr_1332 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_1337;
  assign write_burst_packed_ram_wdata_1337 = _maxi_rdata_sb_0 >> 0;
  assign ram_w8_l262144_id0_0_1_addr = ((write_burst_packed_fsm_25 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_addr_1336 : 'hx;
  assign ram_w8_l262144_id0_0_1_wdata = ((write_burst_packed_fsm_25 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_wdata_1337 : 'hx;
  assign ram_w8_l262144_id0_0_1_wenable = ((write_burst_packed_fsm_25 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  assign ram_w8_l262144_id0_0_1_enable = ((write_burst_packed_fsm_25 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  wire [16-1:0] write_burst_packed_ram_addr_1338;
  assign write_burst_packed_ram_addr_1338 = write_burst_packed_addr_1332 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_1339;
  assign write_burst_packed_ram_wdata_1339 = _maxi_rdata_sb_0 >> 8;
  assign ram_w8_l262144_id0_1_1_addr = ((write_burst_packed_fsm_25 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_addr_1338 : 'hx;
  assign ram_w8_l262144_id0_1_1_wdata = ((write_burst_packed_fsm_25 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_wdata_1339 : 'hx;
  assign ram_w8_l262144_id0_1_1_wenable = ((write_burst_packed_fsm_25 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  assign ram_w8_l262144_id0_1_1_enable = ((write_burst_packed_fsm_25 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  wire [16-1:0] write_burst_packed_ram_addr_1340;
  assign write_burst_packed_ram_addr_1340 = write_burst_packed_addr_1332 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_1341;
  assign write_burst_packed_ram_wdata_1341 = _maxi_rdata_sb_0 >> 16;
  assign ram_w8_l262144_id0_2_1_addr = ((write_burst_packed_fsm_25 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_addr_1340 : 'hx;
  assign ram_w8_l262144_id0_2_1_wdata = ((write_burst_packed_fsm_25 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_wdata_1341 : 'hx;
  assign ram_w8_l262144_id0_2_1_wenable = ((write_burst_packed_fsm_25 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  assign ram_w8_l262144_id0_2_1_enable = ((write_burst_packed_fsm_25 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  wire [16-1:0] write_burst_packed_ram_addr_1342;
  assign write_burst_packed_ram_addr_1342 = write_burst_packed_addr_1332 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_1343;
  assign write_burst_packed_ram_wdata_1343 = _maxi_rdata_sb_0 >> 24;
  assign ram_w8_l262144_id0_3_1_addr = ((write_burst_packed_fsm_25 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_addr_1342 : 'hx;
  assign ram_w8_l262144_id0_3_1_wdata = ((write_burst_packed_fsm_25 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_wdata_1343 : 'hx;
  assign ram_w8_l262144_id0_3_1_wenable = ((write_burst_packed_fsm_25 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  assign ram_w8_l262144_id0_3_1_enable = ((write_burst_packed_fsm_25 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  wire [14-1:0] _dma_read_packed_high_local_size_1344;
  assign _dma_read_packed_high_local_size_1344 = cparam_max_pool_serial_26_act_read_size >> 2;
  wire [2-1:0] _dma_read_packed_low_local_size_1345;
  assign _dma_read_packed_low_local_size_1345 = cparam_max_pool_serial_26_act_read_size & { 2{ 1'd1 } };
  wire [14-1:0] _dma_read_packed_local_packed_size_1346;
  assign _dma_read_packed_local_packed_size_1346 = (_dma_read_packed_low_local_size_1345 > 0)? _dma_read_packed_high_local_size_1344 + 1 : _dma_read_packed_high_local_size_1344;
  wire [32-1:0] mask_addr_shifted_1347;
  assign mask_addr_shifted_1347 = max_pool_serial_26_arg_objaddr_0 + (max_pool_serial_26_act_base_offset + cparam_max_pool_serial_26_act_offset_values_1) + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_1348;
  assign mask_addr_masked_1348 = mask_addr_shifted_1347 << 2;
  reg [32-1:0] max_pool_serial_26_comp_fsm;
  localparam max_pool_serial_26_comp_fsm_init = 0;
  reg [32-1:0] max_pool_serial_26_act_page_comp_offset_buf;
  reg [32-1:0] max_pool_serial_26_out_page_comp_offset_buf;
  reg [32-1:0] max_pool_serial_26_row_count_buf;
  wire max_pool_serial_26_stream_pad_mask_0_0;
  assign max_pool_serial_26_stream_pad_mask_0_0 = (max_pool_serial_26_col_count + 0 < cparam_max_pool_serial_26_pad_col_left) || (max_pool_serial_26_col_count + 0 >= cparam_max_pool_serial_26_act_num_col + cparam_max_pool_serial_26_pad_col_left) || (max_pool_serial_26_row_count_buf + 0 < cparam_max_pool_serial_26_pad_row_top) || (max_pool_serial_26_row_count_buf + 0 >= cparam_max_pool_serial_26_act_num_row + cparam_max_pool_serial_26_pad_row_top);
  wire max_pool_serial_26_stream_pad_mask_0_1;
  assign max_pool_serial_26_stream_pad_mask_0_1 = (max_pool_serial_26_col_count + 1 < cparam_max_pool_serial_26_pad_col_left) || (max_pool_serial_26_col_count + 1 >= cparam_max_pool_serial_26_act_num_col + cparam_max_pool_serial_26_pad_col_left) || (max_pool_serial_26_row_count_buf + 0 < cparam_max_pool_serial_26_pad_row_top) || (max_pool_serial_26_row_count_buf + 0 >= cparam_max_pool_serial_26_act_num_row + cparam_max_pool_serial_26_pad_row_top);
  wire max_pool_serial_26_stream_pad_mask_1_0;
  assign max_pool_serial_26_stream_pad_mask_1_0 = (max_pool_serial_26_col_count + 0 < cparam_max_pool_serial_26_pad_col_left) || (max_pool_serial_26_col_count + 0 >= cparam_max_pool_serial_26_act_num_col + cparam_max_pool_serial_26_pad_col_left) || (max_pool_serial_26_row_count_buf + 1 < cparam_max_pool_serial_26_pad_row_top) || (max_pool_serial_26_row_count_buf + 1 >= cparam_max_pool_serial_26_act_num_row + cparam_max_pool_serial_26_pad_row_top);
  wire max_pool_serial_26_stream_pad_mask_1_1;
  assign max_pool_serial_26_stream_pad_mask_1_1 = (max_pool_serial_26_col_count + 1 < cparam_max_pool_serial_26_pad_col_left) || (max_pool_serial_26_col_count + 1 >= cparam_max_pool_serial_26_act_num_col + cparam_max_pool_serial_26_pad_col_left) || (max_pool_serial_26_row_count_buf + 1 < cparam_max_pool_serial_26_pad_row_top) || (max_pool_serial_26_row_count_buf + 1 >= cparam_max_pool_serial_26_act_num_row + cparam_max_pool_serial_26_pad_row_top);
  reg [4-1:0] max_pool_serial_26_stream_pad_masks;
  wire [3-1:0] stream_max_pool_serial_26_parameter_0_data;
  wire [8-1:0] stream_max_pool_serial_26_source_1_data;
  wire [4-1:0] stream_max_pool_serial_26_parameter_2_data;
  wire [1-1:0] stream_max_pool_serial_26__reduce_reset_data;
  reg __stream_max_pool_serial_26_stream_ivalid_1;
  reg __stream_max_pool_serial_26_stream_ivalid_2;
  reg __stream_max_pool_serial_26_stream_ivalid_3;
  reg __stream_max_pool_serial_26_stream_ivalid_4;
  reg __stream_max_pool_serial_26_stream_ivalid_5;
  reg [32-1:0] _counter_data_897;
  reg [32-1:0] _counter_count_897;
  wire _counter_reset_cond_897;
  assign _counter_reset_cond_897 = stream_max_pool_serial_26__reduce_reset_data;
  wire [32-1:0] _counter_current_count_897;
  assign _counter_current_count_897 = (_counter_reset_cond_897)? 1'sd0 : _counter_count_897;
  wire [8-1:0] _reinterpretcast_src_905;
  assign _reinterpretcast_src_905 = stream_max_pool_serial_26_source_1_data;
  wire signed [8-1:0] _reinterpretcast_data_905;
  assign _reinterpretcast_data_905 = _reinterpretcast_src_905;
  reg [4-1:0] __delay_data_1174__variable_895;
  reg signed [8-1:0] __delay_data_1175_reinterpretcast_905;
  reg [1-1:0] __delay_data_1177__variable_896;
  reg [3-1:0] __delay_data_1180__variable_893;
  reg [1-1:0] _pointer_data_900;
  reg signed [8-1:0] __delay_data_1176__delay_1175_reinterpretcast_905;
  reg [1-1:0] __delay_data_1178__delay_1177__variable_896;
  reg [3-1:0] __delay_data_1181__delay_1180__variable_893;
  reg signed [9-1:0] _cond_data_907;
  reg [1-1:0] __delay_data_1179__delay_1178__delay_1177__variable_896;
  reg [3-1:0] __delay_data_1182__delay_1181__delay_1180__variable_893;
  reg [1-1:0] __variable_wdata_299;
  assign _reduce_max_14__reduce_reset_data = __variable_wdata_299;
  reg signed [8-1:0] __variable_wdata_297;
  assign _reduce_max_14_x_data = __variable_wdata_297;
  reg [32-1:0] __variable_wdata_298;
  assign _reduce_max_14_size_data = __variable_wdata_298;
  assign __reduce_max_14_is_root = ((_stream_max_pool_serial_26_busy)? 0 : 1) && 1;
  assign __reduce_max_14_stream_oready = ((_stream_max_pool_serial_26_busy)? _stream_max_pool_serial_26_stream_oready : 1) && __reduce_max_14_stream_internal_oready;
  assign _stream_max_pool_serial_26_stream_internal_oready = ((_stream_max_pool_serial_26_busy)? __reduce_max_14_stream_internal_oready : 1) && 1;
  wire signed [8-1:0] __substreamoutput_data_909;
  assign __substreamoutput_data_909 = _reduce_max_14_data_data;
  wire [1-1:0] __substreamoutput_data_910;
  assign __substreamoutput_data_910 = _reduce_max_14_valid_data;
  wire signed [8-1:0] _reinterpretcast_src_911;
  assign _reinterpretcast_src_911 = __substreamoutput_data_909;
  wire signed [8-1:0] _reinterpretcast_data_911;
  assign _reinterpretcast_data_911 = _reinterpretcast_src_911;
  wire [1-1:0] stream_max_pool_serial_26_sink_6_data;
  assign stream_max_pool_serial_26_sink_6_data = __substreamoutput_data_910;
  wire signed [8-1:0] stream_max_pool_serial_26_sink_5_data;
  assign stream_max_pool_serial_26_sink_5_data = _reinterpretcast_data_911;
  wire _set_flag_1349;
  assign _set_flag_1349 = max_pool_serial_26_comp_fsm == 4;
  reg [3-1:0] __variable_wdata_893;
  assign stream_max_pool_serial_26_parameter_0_data = __variable_wdata_893;
  wire _set_flag_1350;
  assign _set_flag_1350 = max_pool_serial_26_comp_fsm == 4;
  reg [4-1:0] __variable_wdata_895;
  assign stream_max_pool_serial_26_parameter_2_data = __variable_wdata_895;
  reg [32-1:0] _source_stream_max_pool_serial_26_source_1_pat_cur_offset_0;
  reg [32-1:0] _source_stream_max_pool_serial_26_source_1_pat_cur_offset_1;
  reg [32-1:0] _source_stream_max_pool_serial_26_source_1_pat_cur_offset_2;
  reg [32-1:0] _source_stream_max_pool_serial_26_source_1_pat_cur_offset_3;
  reg [33-1:0] _source_stream_max_pool_serial_26_source_1_pat_size_0;
  reg [33-1:0] _source_stream_max_pool_serial_26_source_1_pat_size_1;
  reg [33-1:0] _source_stream_max_pool_serial_26_source_1_pat_size_2;
  reg [33-1:0] _source_stream_max_pool_serial_26_source_1_pat_size_3;
  reg [32-1:0] _source_stream_max_pool_serial_26_source_1_pat_stride_0;
  reg [32-1:0] _source_stream_max_pool_serial_26_source_1_pat_stride_1;
  reg [32-1:0] _source_stream_max_pool_serial_26_source_1_pat_stride_2;
  reg [32-1:0] _source_stream_max_pool_serial_26_source_1_pat_stride_3;
  reg [33-1:0] _source_stream_max_pool_serial_26_source_1_pat_count_0;
  reg [33-1:0] _source_stream_max_pool_serial_26_source_1_pat_count_1;
  reg [33-1:0] _source_stream_max_pool_serial_26_source_1_pat_count_2;
  reg [33-1:0] _source_stream_max_pool_serial_26_source_1_pat_count_3;
  reg [33-1:0] _source_stream_max_pool_serial_26_source_1_pat_size_buf_0;
  reg [33-1:0] _source_stream_max_pool_serial_26_source_1_pat_size_buf_1;
  reg [33-1:0] _source_stream_max_pool_serial_26_source_1_pat_size_buf_2;
  reg [33-1:0] _source_stream_max_pool_serial_26_source_1_pat_size_buf_3;
  reg [32-1:0] _source_stream_max_pool_serial_26_source_1_pat_stride_buf_0;
  reg [32-1:0] _source_stream_max_pool_serial_26_source_1_pat_stride_buf_1;
  reg [32-1:0] _source_stream_max_pool_serial_26_source_1_pat_stride_buf_2;
  reg [32-1:0] _source_stream_max_pool_serial_26_source_1_pat_stride_buf_3;
  wire _set_flag_1351;
  assign _set_flag_1351 = max_pool_serial_26_comp_fsm == 4;
  wire [2-1:0] read_rtl_bank_1352;
  assign read_rtl_bank_1352 = _stream_max_pool_serial_26_source_1_source_ram_raddr;
  reg [2-1:0] _tmp_1353;
  localparam _tmp_1354 = 1;
  wire [_tmp_1354-1:0] _tmp_1355;
  assign _tmp_1355 = _stream_max_pool_serial_26_stream_oready && _stream_max_pool_serial_26_source_1_source_ram_renable && (_stream_max_pool_serial_26_source_1_source_sel == 1);
  reg [_tmp_1354-1:0] __tmp_1355_1;
  localparam _tmp_1356 = 1;
  wire [_tmp_1356-1:0] _tmp_1357;
  assign _tmp_1357 = _stream_max_pool_serial_26_stream_oready && _stream_max_pool_serial_26_source_1_source_ram_renable && (_stream_max_pool_serial_26_source_1_source_sel == 1);
  reg [_tmp_1356-1:0] __tmp_1357_1;
  localparam _tmp_1358 = 1;
  wire [_tmp_1358-1:0] _tmp_1359;
  assign _tmp_1359 = _stream_max_pool_serial_26_stream_oready && _stream_max_pool_serial_26_source_1_source_ram_renable && (_stream_max_pool_serial_26_source_1_source_sel == 1);
  reg [_tmp_1358-1:0] __tmp_1359_1;
  localparam _tmp_1360 = 1;
  wire [_tmp_1360-1:0] _tmp_1361;
  assign _tmp_1361 = _stream_max_pool_serial_26_stream_oready && _stream_max_pool_serial_26_source_1_source_ram_renable && (_stream_max_pool_serial_26_source_1_source_sel == 1);
  reg [_tmp_1360-1:0] __tmp_1361_1;
  wire signed [8-1:0] read_rtl_rdata_1362;
  wire read_rtl_rvalid_1363;
  assign read_rtl_rdata_1362 = (_tmp_1353 == 0)? ram_w8_l262144_id0_0_0_rdata : 
                               (_tmp_1353 == 1)? ram_w8_l262144_id0_1_0_rdata : 
                               (_tmp_1353 == 2)? ram_w8_l262144_id0_2_0_rdata : 
                               (_tmp_1353 == 3)? ram_w8_l262144_id0_3_0_rdata : 0;
  assign read_rtl_rvalid_1363 = __tmp_1355_1;
  assign _stream_max_pool_serial_26_source_1_source_ram_rdata = (_stream_max_pool_serial_26_source_1_source_sel == 1)? read_rtl_rdata_1362 : 'hx;
  reg [8-1:0] __variable_wdata_894;
  assign stream_max_pool_serial_26_source_1_data = __variable_wdata_894;
  reg [32-1:0] _stream_max_pool_serial_26_source_1_source_pat_fsm_0;
  localparam _stream_max_pool_serial_26_source_1_source_pat_fsm_0_init = 0;
  wire [32-1:0] _stream_max_pool_serial_26_source_1_source_pat_all_offset;
  assign _stream_max_pool_serial_26_source_1_source_pat_all_offset = _stream_max_pool_serial_26_source_1_source_offset_buf + _source_stream_max_pool_serial_26_source_1_pat_cur_offset_0 + _source_stream_max_pool_serial_26_source_1_pat_cur_offset_1 + _source_stream_max_pool_serial_26_source_1_pat_cur_offset_2 + _source_stream_max_pool_serial_26_source_1_pat_cur_offset_3;
  wire _set_flag_1364;
  assign _set_flag_1364 = max_pool_serial_26_comp_fsm == 4;
  reg _tmp_1365;
  reg _tmp_1366;
  reg _tmp_1367;
  reg _tmp_1368;
  reg _tmp_1369;
  reg _tmp_1370;
  reg _tmp_1371;
  localparam _tmp_1372 = 33;
  wire [_tmp_1372-1:0] _tmp_1373;
  assign _tmp_1373 = max_pool_serial_26_stream_out_local + max_pool_serial_26_out_page_comp_offset_buf;
  reg [_tmp_1372-1:0] _tmp_1374;
  reg [_tmp_1372-1:0] _tmp_1375;
  reg [_tmp_1372-1:0] _tmp_1376;
  reg [_tmp_1372-1:0] _tmp_1377;
  reg [_tmp_1372-1:0] _tmp_1378;
  reg [_tmp_1372-1:0] _tmp_1379;
  reg [_tmp_1372-1:0] _tmp_1380;
  reg [10-1:0] _tmp_1381;
  reg [10-1:0] _tmp_1382;
  reg [10-1:0] _tmp_1383;
  reg [10-1:0] _tmp_1384;
  reg [10-1:0] _tmp_1385;
  reg [10-1:0] _tmp_1386;
  reg [10-1:0] _tmp_1387;
  wire [2-1:0] write_rtl_bank_1388;
  assign write_rtl_bank_1388 = _stream_max_pool_serial_26_sink_5_sink_waddr;
  assign ram_w8_l16384_id0_0_0_wdata = (_stream_max_pool_serial_26_stream_oready && _stream_max_pool_serial_26_sink_5_sink_wenable && (_stream_max_pool_serial_26_sink_5_sink_sel == 2) && (write_rtl_bank_1388 == 0))? _stream_max_pool_serial_26_sink_5_sink_wdata : 'hx;
  assign ram_w8_l16384_id0_0_0_wenable = (_stream_max_pool_serial_26_stream_oready && _stream_max_pool_serial_26_sink_5_sink_wenable && (_stream_max_pool_serial_26_sink_5_sink_sel == 2) && (write_rtl_bank_1388 == 0))? 1'd1 : 0;
  assign ram_w8_l16384_id0_1_0_wdata = (_stream_max_pool_serial_26_stream_oready && _stream_max_pool_serial_26_sink_5_sink_wenable && (_stream_max_pool_serial_26_sink_5_sink_sel == 2) && (write_rtl_bank_1388 == 1))? _stream_max_pool_serial_26_sink_5_sink_wdata : 'hx;
  assign ram_w8_l16384_id0_1_0_wenable = (_stream_max_pool_serial_26_stream_oready && _stream_max_pool_serial_26_sink_5_sink_wenable && (_stream_max_pool_serial_26_sink_5_sink_sel == 2) && (write_rtl_bank_1388 == 1))? 1'd1 : 0;
  assign ram_w8_l16384_id0_2_0_wdata = (_stream_max_pool_serial_26_stream_oready && _stream_max_pool_serial_26_sink_5_sink_wenable && (_stream_max_pool_serial_26_sink_5_sink_sel == 2) && (write_rtl_bank_1388 == 2))? _stream_max_pool_serial_26_sink_5_sink_wdata : 'hx;
  assign ram_w8_l16384_id0_2_0_wenable = (_stream_max_pool_serial_26_stream_oready && _stream_max_pool_serial_26_sink_5_sink_wenable && (_stream_max_pool_serial_26_sink_5_sink_sel == 2) && (write_rtl_bank_1388 == 2))? 1'd1 : 0;
  assign ram_w8_l16384_id0_3_0_wdata = (_stream_max_pool_serial_26_stream_oready && _stream_max_pool_serial_26_sink_5_sink_wenable && (_stream_max_pool_serial_26_sink_5_sink_sel == 2) && (write_rtl_bank_1388 == 3))? _stream_max_pool_serial_26_sink_5_sink_wdata : 'hx;
  assign ram_w8_l16384_id0_3_0_wenable = (_stream_max_pool_serial_26_stream_oready && _stream_max_pool_serial_26_sink_5_sink_wenable && (_stream_max_pool_serial_26_sink_5_sink_sel == 2) && (write_rtl_bank_1388 == 3))? 1'd1 : 0;
  reg [32-1:0] _stream_max_pool_serial_26_sink_5_sink_fsm_1;
  localparam _stream_max_pool_serial_26_sink_5_sink_fsm_1_init = 0;
  wire _set_flag_1389;
  assign _set_flag_1389 = max_pool_serial_26_comp_fsm == 5;
  assign _stream_max_pool_serial_26_run_flag = (_set_flag_1389)? 1 : 0;
  reg _tmp_1390;
  reg _tmp_1391;
  reg _tmp_1392;
  reg _tmp_1393;
  reg _tmp_1394;
  reg _tmp_1395;
  reg _tmp_1396;
  reg _tmp_1397;
  reg _tmp_1398;
  reg _tmp_1399;
  assign __reduce_max_14_source_stop = __reduce_max_14_stream_oready && 1'd0;
  reg _tmp_1400;
  reg _tmp_1401;
  reg _tmp_1402;
  assign __reduce_max_14_sink_start = _tmp_1402;
  reg _tmp_1403;
  reg _tmp_1404;
  reg _tmp_1405;
  assign __reduce_max_14_sink_stop = _tmp_1405;
  reg _tmp_1406;
  reg _tmp_1407;
  reg _tmp_1408;
  assign __reduce_max_14_sink_busy = _tmp_1408;
  reg _tmp_1409;
  assign __reduce_max_14_busy = __reduce_max_14_source_busy || __reduce_max_14_sink_busy || __reduce_max_14_busy_reg;
  reg _tmp_1410;
  reg _tmp_1411;
  reg _tmp_1412;
  reg _tmp_1413;
  reg _tmp_1414;
  reg _tmp_1415;
  reg [1-1:0] __variable_wdata_896;
  assign stream_max_pool_serial_26__reduce_reset_data = __variable_wdata_896;
  reg _tmp_1416;
  reg _tmp_1417;
  reg _tmp_1418;
  reg _tmp_1419;
  assign _stream_max_pool_serial_26_source_stop = _stream_max_pool_serial_26_stream_oready && (_stream_max_pool_serial_26_source_1_idle && (_stream_max_pool_serial_26_fsm == 3));
  localparam _tmp_1420 = 1;
  wire [_tmp_1420-1:0] _tmp_1421;
  assign _tmp_1421 = _stream_max_pool_serial_26_source_1_idle && (_stream_max_pool_serial_26_fsm == 3);
  reg [_tmp_1420-1:0] _tmp_1422;
  localparam _tmp_1423 = 1;
  wire [_tmp_1423-1:0] _tmp_1424;
  assign _tmp_1424 = _stream_max_pool_serial_26_source_1_idle && (_stream_max_pool_serial_26_fsm == 3);
  reg [_tmp_1423-1:0] _tmp_1425;
  reg _tmp_1426;
  reg _tmp_1427;
  reg _tmp_1428;
  reg _tmp_1429;
  reg _tmp_1430;
  reg _tmp_1431;
  reg _tmp_1432;
  assign _stream_max_pool_serial_26_sink_start = _tmp_1432;
  reg _tmp_1433;
  reg _tmp_1434;
  reg _tmp_1435;
  reg _tmp_1436;
  reg _tmp_1437;
  reg _tmp_1438;
  reg _tmp_1439;
  assign _stream_max_pool_serial_26_sink_stop = _tmp_1439;
  reg _tmp_1440;
  reg _tmp_1441;
  reg _tmp_1442;
  reg _tmp_1443;
  reg _tmp_1444;
  reg _tmp_1445;
  reg _tmp_1446;
  assign _stream_max_pool_serial_26_sink_busy = _tmp_1446;
  reg _tmp_1447;
  assign _stream_max_pool_serial_26_busy = _stream_max_pool_serial_26_source_busy || _stream_max_pool_serial_26_sink_busy || _stream_max_pool_serial_26_busy_reg;
  wire [13-1:0] _dma_write_packed_high_local_size_1448;
  assign _dma_write_packed_high_local_size_1448 = cparam_max_pool_serial_26_out_write_size >> 2;
  wire [2-1:0] _dma_write_packed_low_local_size_1449;
  assign _dma_write_packed_low_local_size_1449 = cparam_max_pool_serial_26_out_write_size & { 2{ 1'd1 } };
  wire [13-1:0] _dma_write_packed_local_packed_size_1450;
  assign _dma_write_packed_local_packed_size_1450 = (_dma_write_packed_low_local_size_1449 > 0)? _dma_write_packed_high_local_size_1448 + 1 : _dma_write_packed_high_local_size_1448;
  wire [32-1:0] mask_addr_shifted_1451;
  assign mask_addr_shifted_1451 = max_pool_serial_26_objaddr + max_pool_serial_26_out_base_offset + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_1452;
  assign mask_addr_masked_1452 = mask_addr_shifted_1451 << 2;
  reg [32-1:0] read_burst_packed_fsm_26;
  localparam read_burst_packed_fsm_26_init = 0;
  reg [14-1:0] read_burst_packed_addr_1453;
  reg [14-1:0] read_burst_packed_stride_1454;
  reg [33-1:0] read_burst_packed_length_1455;
  reg read_burst_packed_rvalid_1456;
  reg read_burst_packed_rlast_1457;
  wire [12-1:0] read_burst_packed_ram_addr_1458;
  assign read_burst_packed_ram_addr_1458 = read_burst_packed_addr_1453 >> 2;
  localparam _tmp_1459 = 1;
  wire [_tmp_1459-1:0] _tmp_1460;
  assign _tmp_1460 = (read_burst_packed_fsm_26 == 1) && (!read_burst_packed_rvalid_1456 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0));
  reg [_tmp_1459-1:0] __tmp_1460_1;
  wire [8-1:0] read_burst_packed_ram_rdata_1461;
  assign read_burst_packed_ram_rdata_1461 = ram_w8_l16384_id0_0_1_rdata;
  wire [12-1:0] read_burst_packed_ram_addr_1462;
  assign read_burst_packed_ram_addr_1462 = read_burst_packed_addr_1453 >> 2;
  localparam _tmp_1463 = 1;
  wire [_tmp_1463-1:0] _tmp_1464;
  assign _tmp_1464 = (read_burst_packed_fsm_26 == 1) && (!read_burst_packed_rvalid_1456 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0));
  reg [_tmp_1463-1:0] __tmp_1464_1;
  wire [8-1:0] read_burst_packed_ram_rdata_1465;
  assign read_burst_packed_ram_rdata_1465 = ram_w8_l16384_id0_1_1_rdata;
  wire [12-1:0] read_burst_packed_ram_addr_1466;
  assign read_burst_packed_ram_addr_1466 = read_burst_packed_addr_1453 >> 2;
  localparam _tmp_1467 = 1;
  wire [_tmp_1467-1:0] _tmp_1468;
  assign _tmp_1468 = (read_burst_packed_fsm_26 == 1) && (!read_burst_packed_rvalid_1456 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0));
  reg [_tmp_1467-1:0] __tmp_1468_1;
  wire [8-1:0] read_burst_packed_ram_rdata_1469;
  assign read_burst_packed_ram_rdata_1469 = ram_w8_l16384_id0_2_1_rdata;
  wire [12-1:0] read_burst_packed_ram_addr_1470;
  assign read_burst_packed_ram_addr_1470 = read_burst_packed_addr_1453 >> 2;
  localparam _tmp_1471 = 1;
  wire [_tmp_1471-1:0] _tmp_1472;
  assign _tmp_1472 = (read_burst_packed_fsm_26 == 1) && (!read_burst_packed_rvalid_1456 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0));
  reg [_tmp_1471-1:0] __tmp_1472_1;
  wire [8-1:0] read_burst_packed_ram_rdata_1473;
  assign read_burst_packed_ram_rdata_1473 = ram_w8_l16384_id0_3_1_rdata;
  wire [32-1:0] read_burst_packed_rdata_1474;
  assign read_burst_packed_rdata_1474 = { read_burst_packed_ram_rdata_1473, read_burst_packed_ram_rdata_1469, read_burst_packed_ram_rdata_1465, read_burst_packed_ram_rdata_1461 };
  reg _maxi_wdata_cond_1_1;
  reg [32-1:0] avg_pool_serial_52_objaddr;
  reg [32-1:0] avg_pool_serial_52_arg_objaddr_0;
  reg [32-1:0] control_avg_pool_serial_52;
  localparam control_avg_pool_serial_52_init = 0;
  reg _control_avg_pool_serial_52_called;
  wire signed [32-1:0] avg_pool_serial_52_act_base_offset;
  reg signed [32-1:0] avg_pool_serial_52_act_base_offset_row;
  reg signed [32-1:0] avg_pool_serial_52_act_base_offset_bat;
  assign avg_pool_serial_52_act_base_offset = avg_pool_serial_52_act_base_offset_row + avg_pool_serial_52_act_base_offset_bat;
  wire signed [32-1:0] avg_pool_serial_52_out_base_offset;
  reg signed [32-1:0] avg_pool_serial_52_out_base_offset_row;
  reg signed [32-1:0] avg_pool_serial_52_out_base_offset_bat;
  assign avg_pool_serial_52_out_base_offset = avg_pool_serial_52_out_base_offset_row + avg_pool_serial_52_out_base_offset_bat;
  reg [32-1:0] avg_pool_serial_52_col_count;
  reg [32-1:0] avg_pool_serial_52_row_count;
  reg [32-1:0] avg_pool_serial_52_bat_count;
  reg [32-1:0] avg_pool_serial_52_prev_row_count;
  reg [32-1:0] avg_pool_serial_52_prev_bat_count;
  reg [32-1:0] avg_pool_serial_52_stream_act_local;
  reg [32-1:0] avg_pool_serial_52_stream_out_local;
  reg avg_pool_serial_52_act_page;
  reg [32-1:0] avg_pool_serial_52_act_page_comp_offset;
  reg [32-1:0] avg_pool_serial_52_act_page_dma_offset;
  reg avg_pool_serial_52_out_page;
  reg [32-1:0] avg_pool_serial_52_out_page_comp_offset;
  reg [32-1:0] avg_pool_serial_52_out_page_dma_offset;
  reg avg_pool_serial_52_skip_read_act;
  reg avg_pool_serial_52_skip_comp;
  reg avg_pool_serial_52_skip_write_out;
  reg [32-1:0] avg_pool_serial_52_comp_count;
  reg [32-1:0] avg_pool_serial_52_out_count;
  wire avg_pool_serial_52_dma_pad_mask_0;
  assign avg_pool_serial_52_dma_pad_mask_0 = (avg_pool_serial_52_row_count + 0 < cparam_avg_pool_serial_52_pad_row_top) || (avg_pool_serial_52_row_count + 0 >= cparam_avg_pool_serial_52_act_num_row + cparam_avg_pool_serial_52_pad_row_top);
  wire [12-1:0] _dma_read_packed_high_local_size_1475;
  assign _dma_read_packed_high_local_size_1475 = cparam_avg_pool_serial_52_act_read_size >> 2;
  wire [2-1:0] _dma_read_packed_low_local_size_1476;
  assign _dma_read_packed_low_local_size_1476 = cparam_avg_pool_serial_52_act_read_size & { 2{ 1'd1 } };
  wire [12-1:0] _dma_read_packed_local_packed_size_1477;
  assign _dma_read_packed_local_packed_size_1477 = (_dma_read_packed_low_local_size_1476 > 0)? _dma_read_packed_high_local_size_1475 + 1 : _dma_read_packed_high_local_size_1475;
  wire [32-1:0] mask_addr_shifted_1478;
  assign mask_addr_shifted_1478 = avg_pool_serial_52_arg_objaddr_0 + (avg_pool_serial_52_act_base_offset + cparam_avg_pool_serial_52_act_offset_values_0) + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_1479;
  assign mask_addr_masked_1479 = mask_addr_shifted_1478 << 2;
  reg [32-1:0] write_burst_packed_fsm_27;
  localparam write_burst_packed_fsm_27_init = 0;
  reg [14-1:0] write_burst_packed_addr_1480;
  reg [14-1:0] write_burst_packed_stride_1481;
  reg [33-1:0] write_burst_packed_length_1482;
  reg write_burst_packed_done_1483;
  wire [12-1:0] write_burst_packed_ram_addr_1484;
  assign write_burst_packed_ram_addr_1484 = write_burst_packed_addr_1480 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_1485;
  assign write_burst_packed_ram_wdata_1485 = _maxi_rdata_sb_0 >> 0;
  assign ram_w8_l16384_id0_0_1_addr = ((write_burst_packed_fsm_27 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_addr_1484 : 
                                      ((read_burst_packed_fsm_26 == 1) && (!read_burst_packed_rvalid_1456 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)))? read_burst_packed_ram_addr_1458 : 
                                      ((write_burst_packed_fsm_12 == 1) && write_burst_block_ram_wvalid_243)? write_burst_packed_ram_addr_249 : 'hx;
  assign ram_w8_l16384_id0_0_1_wdata = ((write_burst_packed_fsm_27 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_wdata_1485 : 
                                       ((write_burst_packed_fsm_12 == 1) && write_burst_block_ram_wvalid_243)? write_burst_packed_ram_wdata_250 : 'hx;
  assign ram_w8_l16384_id0_0_1_wenable = ((write_burst_packed_fsm_27 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 
                                         ((write_burst_packed_fsm_12 == 1) && write_burst_block_ram_wvalid_243)? 1'd1 : 0;
  assign ram_w8_l16384_id0_0_1_enable = ((write_burst_packed_fsm_27 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 
                                        ((read_burst_packed_fsm_26 == 1) && (!read_burst_packed_rvalid_1456 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)))? 1'd1 : 
                                        ((write_burst_packed_fsm_12 == 1) && write_burst_block_ram_wvalid_243)? 1'd1 : 0;
  wire [12-1:0] write_burst_packed_ram_addr_1486;
  assign write_burst_packed_ram_addr_1486 = write_burst_packed_addr_1480 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_1487;
  assign write_burst_packed_ram_wdata_1487 = _maxi_rdata_sb_0 >> 8;
  assign ram_w8_l16384_id0_1_1_addr = ((write_burst_packed_fsm_27 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_addr_1486 : 
                                      ((read_burst_packed_fsm_26 == 1) && (!read_burst_packed_rvalid_1456 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)))? read_burst_packed_ram_addr_1462 : 
                                      ((write_burst_packed_fsm_12 == 1) && write_burst_block_ram_wvalid_243)? write_burst_packed_ram_addr_251 : 'hx;
  assign ram_w8_l16384_id0_1_1_wdata = ((write_burst_packed_fsm_27 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_wdata_1487 : 
                                       ((write_burst_packed_fsm_12 == 1) && write_burst_block_ram_wvalid_243)? write_burst_packed_ram_wdata_252 : 'hx;
  assign ram_w8_l16384_id0_1_1_wenable = ((write_burst_packed_fsm_27 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 
                                         ((write_burst_packed_fsm_12 == 1) && write_burst_block_ram_wvalid_243)? 1'd1 : 0;
  assign ram_w8_l16384_id0_1_1_enable = ((write_burst_packed_fsm_27 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 
                                        ((read_burst_packed_fsm_26 == 1) && (!read_burst_packed_rvalid_1456 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)))? 1'd1 : 
                                        ((write_burst_packed_fsm_12 == 1) && write_burst_block_ram_wvalid_243)? 1'd1 : 0;
  wire [12-1:0] write_burst_packed_ram_addr_1488;
  assign write_burst_packed_ram_addr_1488 = write_burst_packed_addr_1480 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_1489;
  assign write_burst_packed_ram_wdata_1489 = _maxi_rdata_sb_0 >> 16;
  assign ram_w8_l16384_id0_2_1_addr = ((write_burst_packed_fsm_27 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_addr_1488 : 
                                      ((read_burst_packed_fsm_26 == 1) && (!read_burst_packed_rvalid_1456 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)))? read_burst_packed_ram_addr_1466 : 
                                      ((write_burst_packed_fsm_12 == 1) && write_burst_block_ram_wvalid_243)? write_burst_packed_ram_addr_253 : 'hx;
  assign ram_w8_l16384_id0_2_1_wdata = ((write_burst_packed_fsm_27 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_wdata_1489 : 
                                       ((write_burst_packed_fsm_12 == 1) && write_burst_block_ram_wvalid_243)? write_burst_packed_ram_wdata_254 : 'hx;
  assign ram_w8_l16384_id0_2_1_wenable = ((write_burst_packed_fsm_27 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 
                                         ((write_burst_packed_fsm_12 == 1) && write_burst_block_ram_wvalid_243)? 1'd1 : 0;
  assign ram_w8_l16384_id0_2_1_enable = ((write_burst_packed_fsm_27 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 
                                        ((read_burst_packed_fsm_26 == 1) && (!read_burst_packed_rvalid_1456 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)))? 1'd1 : 
                                        ((write_burst_packed_fsm_12 == 1) && write_burst_block_ram_wvalid_243)? 1'd1 : 0;
  wire [12-1:0] write_burst_packed_ram_addr_1490;
  assign write_burst_packed_ram_addr_1490 = write_burst_packed_addr_1480 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_1491;
  assign write_burst_packed_ram_wdata_1491 = _maxi_rdata_sb_0 >> 24;
  assign ram_w8_l16384_id0_3_1_addr = ((write_burst_packed_fsm_27 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_addr_1490 : 
                                      ((read_burst_packed_fsm_26 == 1) && (!read_burst_packed_rvalid_1456 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)))? read_burst_packed_ram_addr_1470 : 
                                      ((write_burst_packed_fsm_12 == 1) && write_burst_block_ram_wvalid_243)? write_burst_packed_ram_addr_255 : 'hx;
  assign ram_w8_l16384_id0_3_1_wdata = ((write_burst_packed_fsm_27 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_wdata_1491 : 
                                       ((write_burst_packed_fsm_12 == 1) && write_burst_block_ram_wvalid_243)? write_burst_packed_ram_wdata_256 : 'hx;
  assign ram_w8_l16384_id0_3_1_wenable = ((write_burst_packed_fsm_27 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 
                                         ((write_burst_packed_fsm_12 == 1) && write_burst_block_ram_wvalid_243)? 1'd1 : 0;
  assign ram_w8_l16384_id0_3_1_enable = ((write_burst_packed_fsm_27 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 
                                        ((read_burst_packed_fsm_26 == 1) && (!read_burst_packed_rvalid_1456 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)))? 1'd1 : 
                                        ((write_burst_packed_fsm_12 == 1) && write_burst_block_ram_wvalid_243)? 1'd1 : 0;
  reg [32-1:0] avg_pool_serial_52_comp_fsm;
  localparam avg_pool_serial_52_comp_fsm_init = 0;
  reg [32-1:0] avg_pool_serial_52_act_page_comp_offset_buf;
  reg [32-1:0] avg_pool_serial_52_out_page_comp_offset_buf;
  reg [32-1:0] avg_pool_serial_52_row_count_buf;
  wire avg_pool_serial_52_stream_pad_mask_0_0;
  assign avg_pool_serial_52_stream_pad_mask_0_0 = (avg_pool_serial_52_col_count + 0 < cparam_avg_pool_serial_52_pad_col_left) || (avg_pool_serial_52_col_count + 0 >= cparam_avg_pool_serial_52_act_num_col + cparam_avg_pool_serial_52_pad_col_left) || (avg_pool_serial_52_row_count_buf + 0 < cparam_avg_pool_serial_52_pad_row_top) || (avg_pool_serial_52_row_count_buf + 0 >= cparam_avg_pool_serial_52_act_num_row + cparam_avg_pool_serial_52_pad_row_top);
  reg [1-1:0] avg_pool_serial_52_stream_pad_masks;
  wire [1-1:0] stream_avg_pool_serial_52_parameter_0_data;
  wire [8-1:0] stream_avg_pool_serial_52_source_1_data;
  wire [1-1:0] stream_avg_pool_serial_52_parameter_2_data;
  wire [1-1:0] stream_avg_pool_serial_52__reduce_reset_data;
  reg __stream_avg_pool_serial_52_stream_ivalid_1;
  reg __stream_avg_pool_serial_52_stream_ivalid_2;
  reg __stream_avg_pool_serial_52_stream_ivalid_3;
  reg __stream_avg_pool_serial_52_stream_ivalid_4;
  reg __stream_avg_pool_serial_52_stream_ivalid_5;
  reg __stream_avg_pool_serial_52_stream_ivalid_6;
  reg [32-1:0] _counter_data_916;
  reg [32-1:0] _counter_count_916;
  wire _counter_reset_cond_916;
  assign _counter_reset_cond_916 = stream_avg_pool_serial_52__reduce_reset_data;
  wire [32-1:0] _counter_current_count_916;
  assign _counter_current_count_916 = (_counter_reset_cond_916)? 1'sd0 : _counter_count_916;
  wire [8-1:0] _reinterpretcast_src_924;
  assign _reinterpretcast_src_924 = stream_avg_pool_serial_52_source_1_data;
  wire signed [8-1:0] _reinterpretcast_data_924;
  assign _reinterpretcast_data_924 = _reinterpretcast_src_924;
  reg [1-1:0] __delay_data_1183__variable_914;
  reg signed [8-1:0] __delay_data_1184_reinterpretcast_924;
  reg [1-1:0] __delay_data_1186__variable_915;
  reg [1-1:0] __delay_data_1189__variable_912;
  reg [1-1:0] _pointer_data_919;
  reg signed [8-1:0] __delay_data_1185__delay_1184_reinterpretcast_924;
  reg [1-1:0] __delay_data_1187__delay_1186__variable_915;
  reg [1-1:0] __delay_data_1190__delay_1189__variable_912;
  reg signed [8-1:0] _cond_data_926;
  reg [1-1:0] __delay_data_1188__delay_1187__delay_1186__variable_915;
  reg [1-1:0] __delay_data_1191__delay_1190__delay_1189__variable_912;
  reg [1-1:0] __variable_wdata_3;
  assign acc_0__reduce_reset_data = __variable_wdata_3;
  reg signed [32-1:0] __variable_wdata_0;
  assign acc_0_x_data = __variable_wdata_0;
  reg [32-1:0] __variable_wdata_2;
  assign acc_0_size_data = __variable_wdata_2;
  reg [6-1:0] __variable_wdata_1;
  assign acc_0_rshift_data = __variable_wdata_1;
  assign _acc_0_is_root = ((_stream_avg_pool_serial_52_busy)? 0 : 1) && 1;
  assign _acc_0_stream_oready = ((_stream_avg_pool_serial_52_busy)? _stream_avg_pool_serial_52_stream_oready : 1) && _acc_0_stream_internal_oready;
  assign _stream_avg_pool_serial_52_stream_internal_oready = ((_stream_avg_pool_serial_52_busy)? _acc_0_stream_internal_oready : 1) && 1;
  wire signed [32-1:0] __substreamoutput_data_932;
  assign __substreamoutput_data_932 = acc_0_sum_data;
  wire [1-1:0] __substreamoutput_data_933;
  assign __substreamoutput_data_933 = acc_0_valid_data;
  wire signed [32-1:0] _reinterpretcast_src_935;
  assign _reinterpretcast_src_935 = __substreamoutput_data_932;
  wire signed [8-1:0] _reinterpretcast_data_935;
  assign _reinterpretcast_data_935 = _reinterpretcast_src_935;
  wire [1-1:0] stream_avg_pool_serial_52_sink_6_data;
  assign stream_avg_pool_serial_52_sink_6_data = __substreamoutput_data_933;
  wire signed [8-1:0] stream_avg_pool_serial_52_sink_5_data;
  assign stream_avg_pool_serial_52_sink_5_data = _reinterpretcast_data_935;
  wire _set_flag_1492;
  assign _set_flag_1492 = avg_pool_serial_52_comp_fsm == 4;
  reg [1-1:0] __variable_wdata_912;
  assign stream_avg_pool_serial_52_parameter_0_data = __variable_wdata_912;
  wire _set_flag_1493;
  assign _set_flag_1493 = avg_pool_serial_52_comp_fsm == 4;
  reg [1-1:0] __variable_wdata_914;
  assign stream_avg_pool_serial_52_parameter_2_data = __variable_wdata_914;
  reg [32-1:0] _source_stream_avg_pool_serial_52_source_1_pat_cur_offset_0;
  reg [32-1:0] _source_stream_avg_pool_serial_52_source_1_pat_cur_offset_1;
  reg [32-1:0] _source_stream_avg_pool_serial_52_source_1_pat_cur_offset_2;
  reg [32-1:0] _source_stream_avg_pool_serial_52_source_1_pat_cur_offset_3;
  reg [33-1:0] _source_stream_avg_pool_serial_52_source_1_pat_size_0;
  reg [33-1:0] _source_stream_avg_pool_serial_52_source_1_pat_size_1;
  reg [33-1:0] _source_stream_avg_pool_serial_52_source_1_pat_size_2;
  reg [33-1:0] _source_stream_avg_pool_serial_52_source_1_pat_size_3;
  reg [32-1:0] _source_stream_avg_pool_serial_52_source_1_pat_stride_0;
  reg [32-1:0] _source_stream_avg_pool_serial_52_source_1_pat_stride_1;
  reg [32-1:0] _source_stream_avg_pool_serial_52_source_1_pat_stride_2;
  reg [32-1:0] _source_stream_avg_pool_serial_52_source_1_pat_stride_3;
  reg [33-1:0] _source_stream_avg_pool_serial_52_source_1_pat_count_0;
  reg [33-1:0] _source_stream_avg_pool_serial_52_source_1_pat_count_1;
  reg [33-1:0] _source_stream_avg_pool_serial_52_source_1_pat_count_2;
  reg [33-1:0] _source_stream_avg_pool_serial_52_source_1_pat_count_3;
  reg [33-1:0] _source_stream_avg_pool_serial_52_source_1_pat_size_buf_0;
  reg [33-1:0] _source_stream_avg_pool_serial_52_source_1_pat_size_buf_1;
  reg [33-1:0] _source_stream_avg_pool_serial_52_source_1_pat_size_buf_2;
  reg [33-1:0] _source_stream_avg_pool_serial_52_source_1_pat_size_buf_3;
  reg [32-1:0] _source_stream_avg_pool_serial_52_source_1_pat_stride_buf_0;
  reg [32-1:0] _source_stream_avg_pool_serial_52_source_1_pat_stride_buf_1;
  reg [32-1:0] _source_stream_avg_pool_serial_52_source_1_pat_stride_buf_2;
  reg [32-1:0] _source_stream_avg_pool_serial_52_source_1_pat_stride_buf_3;
  wire _set_flag_1494;
  assign _set_flag_1494 = avg_pool_serial_52_comp_fsm == 4;
  wire [2-1:0] read_rtl_bank_1495;
  assign read_rtl_bank_1495 = _stream_avg_pool_serial_52_source_1_source_ram_raddr;
  reg [2-1:0] _tmp_1496;
  assign ram_w8_l16384_id0_0_0_addr = (_stream_avg_pool_serial_52_stream_oready && _stream_avg_pool_serial_52_source_1_source_ram_renable && (_stream_avg_pool_serial_52_source_1_source_sel == 1))? _stream_avg_pool_serial_52_source_1_source_ram_raddr >> 2 : 
                                      (_stream_max_pool_serial_26_stream_oready && _stream_max_pool_serial_26_sink_5_sink_wenable && (_stream_max_pool_serial_26_sink_5_sink_sel == 2) && (write_rtl_bank_1388 == 0))? _stream_max_pool_serial_26_sink_5_sink_waddr >> 2 : 
                                      (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_20_source_ram_renable && (_stream_conv2d_24_source_20_source_sel == 3))? _stream_conv2d_24_source_20_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l16384_id0_0_0_enable = (_stream_avg_pool_serial_52_stream_oready && _stream_avg_pool_serial_52_source_1_source_ram_renable && (_stream_avg_pool_serial_52_source_1_source_sel == 1))? 1'd1 : 
                                        (_stream_max_pool_serial_26_stream_oready && _stream_max_pool_serial_26_sink_5_sink_wenable && (_stream_max_pool_serial_26_sink_5_sink_sel == 2) && (write_rtl_bank_1388 == 0))? 1'd1 : 
                                        (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_20_source_ram_renable && (_stream_conv2d_24_source_20_source_sel == 3))? 1'd1 : 0;
  localparam _tmp_1497 = 1;
  wire [_tmp_1497-1:0] _tmp_1498;
  assign _tmp_1498 = _stream_avg_pool_serial_52_stream_oready && _stream_avg_pool_serial_52_source_1_source_ram_renable && (_stream_avg_pool_serial_52_source_1_source_sel == 1);
  reg [_tmp_1497-1:0] __tmp_1498_1;
  assign ram_w8_l16384_id0_1_0_addr = (_stream_avg_pool_serial_52_stream_oready && _stream_avg_pool_serial_52_source_1_source_ram_renable && (_stream_avg_pool_serial_52_source_1_source_sel == 1))? _stream_avg_pool_serial_52_source_1_source_ram_raddr >> 2 : 
                                      (_stream_max_pool_serial_26_stream_oready && _stream_max_pool_serial_26_sink_5_sink_wenable && (_stream_max_pool_serial_26_sink_5_sink_sel == 2) && (write_rtl_bank_1388 == 1))? _stream_max_pool_serial_26_sink_5_sink_waddr >> 2 : 
                                      (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_20_source_ram_renable && (_stream_conv2d_24_source_20_source_sel == 3))? _stream_conv2d_24_source_20_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l16384_id0_1_0_enable = (_stream_avg_pool_serial_52_stream_oready && _stream_avg_pool_serial_52_source_1_source_ram_renable && (_stream_avg_pool_serial_52_source_1_source_sel == 1))? 1'd1 : 
                                        (_stream_max_pool_serial_26_stream_oready && _stream_max_pool_serial_26_sink_5_sink_wenable && (_stream_max_pool_serial_26_sink_5_sink_sel == 2) && (write_rtl_bank_1388 == 1))? 1'd1 : 
                                        (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_20_source_ram_renable && (_stream_conv2d_24_source_20_source_sel == 3))? 1'd1 : 0;
  localparam _tmp_1499 = 1;
  wire [_tmp_1499-1:0] _tmp_1500;
  assign _tmp_1500 = _stream_avg_pool_serial_52_stream_oready && _stream_avg_pool_serial_52_source_1_source_ram_renable && (_stream_avg_pool_serial_52_source_1_source_sel == 1);
  reg [_tmp_1499-1:0] __tmp_1500_1;
  assign ram_w8_l16384_id0_2_0_addr = (_stream_avg_pool_serial_52_stream_oready && _stream_avg_pool_serial_52_source_1_source_ram_renable && (_stream_avg_pool_serial_52_source_1_source_sel == 1))? _stream_avg_pool_serial_52_source_1_source_ram_raddr >> 2 : 
                                      (_stream_max_pool_serial_26_stream_oready && _stream_max_pool_serial_26_sink_5_sink_wenable && (_stream_max_pool_serial_26_sink_5_sink_sel == 2) && (write_rtl_bank_1388 == 2))? _stream_max_pool_serial_26_sink_5_sink_waddr >> 2 : 
                                      (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_20_source_ram_renable && (_stream_conv2d_24_source_20_source_sel == 3))? _stream_conv2d_24_source_20_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l16384_id0_2_0_enable = (_stream_avg_pool_serial_52_stream_oready && _stream_avg_pool_serial_52_source_1_source_ram_renable && (_stream_avg_pool_serial_52_source_1_source_sel == 1))? 1'd1 : 
                                        (_stream_max_pool_serial_26_stream_oready && _stream_max_pool_serial_26_sink_5_sink_wenable && (_stream_max_pool_serial_26_sink_5_sink_sel == 2) && (write_rtl_bank_1388 == 2))? 1'd1 : 
                                        (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_20_source_ram_renable && (_stream_conv2d_24_source_20_source_sel == 3))? 1'd1 : 0;
  localparam _tmp_1501 = 1;
  wire [_tmp_1501-1:0] _tmp_1502;
  assign _tmp_1502 = _stream_avg_pool_serial_52_stream_oready && _stream_avg_pool_serial_52_source_1_source_ram_renable && (_stream_avg_pool_serial_52_source_1_source_sel == 1);
  reg [_tmp_1501-1:0] __tmp_1502_1;
  assign ram_w8_l16384_id0_3_0_addr = (_stream_avg_pool_serial_52_stream_oready && _stream_avg_pool_serial_52_source_1_source_ram_renable && (_stream_avg_pool_serial_52_source_1_source_sel == 1))? _stream_avg_pool_serial_52_source_1_source_ram_raddr >> 2 : 
                                      (_stream_max_pool_serial_26_stream_oready && _stream_max_pool_serial_26_sink_5_sink_wenable && (_stream_max_pool_serial_26_sink_5_sink_sel == 2) && (write_rtl_bank_1388 == 3))? _stream_max_pool_serial_26_sink_5_sink_waddr >> 2 : 
                                      (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_20_source_ram_renable && (_stream_conv2d_24_source_20_source_sel == 3))? _stream_conv2d_24_source_20_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l16384_id0_3_0_enable = (_stream_avg_pool_serial_52_stream_oready && _stream_avg_pool_serial_52_source_1_source_ram_renable && (_stream_avg_pool_serial_52_source_1_source_sel == 1))? 1'd1 : 
                                        (_stream_max_pool_serial_26_stream_oready && _stream_max_pool_serial_26_sink_5_sink_wenable && (_stream_max_pool_serial_26_sink_5_sink_sel == 2) && (write_rtl_bank_1388 == 3))? 1'd1 : 
                                        (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_20_source_ram_renable && (_stream_conv2d_24_source_20_source_sel == 3))? 1'd1 : 0;
  localparam _tmp_1503 = 1;
  wire [_tmp_1503-1:0] _tmp_1504;
  assign _tmp_1504 = _stream_avg_pool_serial_52_stream_oready && _stream_avg_pool_serial_52_source_1_source_ram_renable && (_stream_avg_pool_serial_52_source_1_source_sel == 1);
  reg [_tmp_1503-1:0] __tmp_1504_1;
  wire signed [8-1:0] read_rtl_rdata_1505;
  wire read_rtl_rvalid_1506;
  assign read_rtl_rdata_1505 = (_tmp_1496 == 0)? ram_w8_l16384_id0_0_0_rdata : 
                               (_tmp_1496 == 1)? ram_w8_l16384_id0_1_0_rdata : 
                               (_tmp_1496 == 2)? ram_w8_l16384_id0_2_0_rdata : 
                               (_tmp_1496 == 3)? ram_w8_l16384_id0_3_0_rdata : 0;
  assign read_rtl_rvalid_1506 = __tmp_1498_1;
  assign _stream_avg_pool_serial_52_source_1_source_ram_rdata = (_stream_avg_pool_serial_52_source_1_source_sel == 1)? read_rtl_rdata_1505 : 'hx;
  reg [8-1:0] __variable_wdata_913;
  assign stream_avg_pool_serial_52_source_1_data = __variable_wdata_913;
  reg [32-1:0] _stream_avg_pool_serial_52_source_1_source_pat_fsm_0;
  localparam _stream_avg_pool_serial_52_source_1_source_pat_fsm_0_init = 0;
  wire [32-1:0] _stream_avg_pool_serial_52_source_1_source_pat_all_offset;
  assign _stream_avg_pool_serial_52_source_1_source_pat_all_offset = _stream_avg_pool_serial_52_source_1_source_offset_buf + _source_stream_avg_pool_serial_52_source_1_pat_cur_offset_0 + _source_stream_avg_pool_serial_52_source_1_pat_cur_offset_1 + _source_stream_avg_pool_serial_52_source_1_pat_cur_offset_2 + _source_stream_avg_pool_serial_52_source_1_pat_cur_offset_3;
  wire _set_flag_1507;
  assign _set_flag_1507 = avg_pool_serial_52_comp_fsm == 4;
  reg _tmp_1508;
  reg _tmp_1509;
  reg _tmp_1510;
  reg _tmp_1511;
  reg _tmp_1512;
  reg _tmp_1513;
  reg _tmp_1514;
  reg _tmp_1515;
  localparam _tmp_1516 = 33;
  wire [_tmp_1516-1:0] _tmp_1517;
  assign _tmp_1517 = avg_pool_serial_52_stream_out_local + avg_pool_serial_52_out_page_comp_offset_buf;
  reg [_tmp_1516-1:0] _tmp_1518;
  reg [_tmp_1516-1:0] _tmp_1519;
  reg [_tmp_1516-1:0] _tmp_1520;
  reg [_tmp_1516-1:0] _tmp_1521;
  reg [_tmp_1516-1:0] _tmp_1522;
  reg [_tmp_1516-1:0] _tmp_1523;
  reg [_tmp_1516-1:0] _tmp_1524;
  reg [_tmp_1516-1:0] _tmp_1525;
  reg [10-1:0] _tmp_1526;
  reg [10-1:0] _tmp_1527;
  reg [10-1:0] _tmp_1528;
  reg [10-1:0] _tmp_1529;
  reg [10-1:0] _tmp_1530;
  reg [10-1:0] _tmp_1531;
  reg [10-1:0] _tmp_1532;
  reg [10-1:0] _tmp_1533;
  wire [2-1:0] write_rtl_bank_1534;
  assign write_rtl_bank_1534 = _stream_avg_pool_serial_52_sink_5_sink_waddr;
  assign ram_w8_l16384_id1_0_0_addr = (_stream_avg_pool_serial_52_stream_oready && _stream_avg_pool_serial_52_sink_5_sink_wenable && (_stream_avg_pool_serial_52_sink_5_sink_sel == 2) && (write_rtl_bank_1534 == 0))? _stream_avg_pool_serial_52_sink_5_sink_waddr >> 2 : 
                                      (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_21_source_ram_renable && (_stream_conv2d_24_source_21_source_sel == 4))? _stream_conv2d_24_source_21_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l16384_id1_0_0_wdata = (_stream_avg_pool_serial_52_stream_oready && _stream_avg_pool_serial_52_sink_5_sink_wenable && (_stream_avg_pool_serial_52_sink_5_sink_sel == 2) && (write_rtl_bank_1534 == 0))? _stream_avg_pool_serial_52_sink_5_sink_wdata : 'hx;
  assign ram_w8_l16384_id1_0_0_wenable = (_stream_avg_pool_serial_52_stream_oready && _stream_avg_pool_serial_52_sink_5_sink_wenable && (_stream_avg_pool_serial_52_sink_5_sink_sel == 2) && (write_rtl_bank_1534 == 0))? 1'd1 : 0;
  assign ram_w8_l16384_id1_0_0_enable = (_stream_avg_pool_serial_52_stream_oready && _stream_avg_pool_serial_52_sink_5_sink_wenable && (_stream_avg_pool_serial_52_sink_5_sink_sel == 2) && (write_rtl_bank_1534 == 0))? 1'd1 : 
                                        (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_21_source_ram_renable && (_stream_conv2d_24_source_21_source_sel == 4))? 1'd1 : 0;
  assign ram_w8_l16384_id1_1_0_addr = (_stream_avg_pool_serial_52_stream_oready && _stream_avg_pool_serial_52_sink_5_sink_wenable && (_stream_avg_pool_serial_52_sink_5_sink_sel == 2) && (write_rtl_bank_1534 == 1))? _stream_avg_pool_serial_52_sink_5_sink_waddr >> 2 : 
                                      (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_21_source_ram_renable && (_stream_conv2d_24_source_21_source_sel == 4))? _stream_conv2d_24_source_21_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l16384_id1_1_0_wdata = (_stream_avg_pool_serial_52_stream_oready && _stream_avg_pool_serial_52_sink_5_sink_wenable && (_stream_avg_pool_serial_52_sink_5_sink_sel == 2) && (write_rtl_bank_1534 == 1))? _stream_avg_pool_serial_52_sink_5_sink_wdata : 'hx;
  assign ram_w8_l16384_id1_1_0_wenable = (_stream_avg_pool_serial_52_stream_oready && _stream_avg_pool_serial_52_sink_5_sink_wenable && (_stream_avg_pool_serial_52_sink_5_sink_sel == 2) && (write_rtl_bank_1534 == 1))? 1'd1 : 0;
  assign ram_w8_l16384_id1_1_0_enable = (_stream_avg_pool_serial_52_stream_oready && _stream_avg_pool_serial_52_sink_5_sink_wenable && (_stream_avg_pool_serial_52_sink_5_sink_sel == 2) && (write_rtl_bank_1534 == 1))? 1'd1 : 
                                        (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_21_source_ram_renable && (_stream_conv2d_24_source_21_source_sel == 4))? 1'd1 : 0;
  assign ram_w8_l16384_id1_2_0_addr = (_stream_avg_pool_serial_52_stream_oready && _stream_avg_pool_serial_52_sink_5_sink_wenable && (_stream_avg_pool_serial_52_sink_5_sink_sel == 2) && (write_rtl_bank_1534 == 2))? _stream_avg_pool_serial_52_sink_5_sink_waddr >> 2 : 
                                      (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_21_source_ram_renable && (_stream_conv2d_24_source_21_source_sel == 4))? _stream_conv2d_24_source_21_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l16384_id1_2_0_wdata = (_stream_avg_pool_serial_52_stream_oready && _stream_avg_pool_serial_52_sink_5_sink_wenable && (_stream_avg_pool_serial_52_sink_5_sink_sel == 2) && (write_rtl_bank_1534 == 2))? _stream_avg_pool_serial_52_sink_5_sink_wdata : 'hx;
  assign ram_w8_l16384_id1_2_0_wenable = (_stream_avg_pool_serial_52_stream_oready && _stream_avg_pool_serial_52_sink_5_sink_wenable && (_stream_avg_pool_serial_52_sink_5_sink_sel == 2) && (write_rtl_bank_1534 == 2))? 1'd1 : 0;
  assign ram_w8_l16384_id1_2_0_enable = (_stream_avg_pool_serial_52_stream_oready && _stream_avg_pool_serial_52_sink_5_sink_wenable && (_stream_avg_pool_serial_52_sink_5_sink_sel == 2) && (write_rtl_bank_1534 == 2))? 1'd1 : 
                                        (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_21_source_ram_renable && (_stream_conv2d_24_source_21_source_sel == 4))? 1'd1 : 0;
  assign ram_w8_l16384_id1_3_0_addr = (_stream_avg_pool_serial_52_stream_oready && _stream_avg_pool_serial_52_sink_5_sink_wenable && (_stream_avg_pool_serial_52_sink_5_sink_sel == 2) && (write_rtl_bank_1534 == 3))? _stream_avg_pool_serial_52_sink_5_sink_waddr >> 2 : 
                                      (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_21_source_ram_renable && (_stream_conv2d_24_source_21_source_sel == 4))? _stream_conv2d_24_source_21_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l16384_id1_3_0_wdata = (_stream_avg_pool_serial_52_stream_oready && _stream_avg_pool_serial_52_sink_5_sink_wenable && (_stream_avg_pool_serial_52_sink_5_sink_sel == 2) && (write_rtl_bank_1534 == 3))? _stream_avg_pool_serial_52_sink_5_sink_wdata : 'hx;
  assign ram_w8_l16384_id1_3_0_wenable = (_stream_avg_pool_serial_52_stream_oready && _stream_avg_pool_serial_52_sink_5_sink_wenable && (_stream_avg_pool_serial_52_sink_5_sink_sel == 2) && (write_rtl_bank_1534 == 3))? 1'd1 : 0;
  assign ram_w8_l16384_id1_3_0_enable = (_stream_avg_pool_serial_52_stream_oready && _stream_avg_pool_serial_52_sink_5_sink_wenable && (_stream_avg_pool_serial_52_sink_5_sink_sel == 2) && (write_rtl_bank_1534 == 3))? 1'd1 : 
                                        (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_21_source_ram_renable && (_stream_conv2d_24_source_21_source_sel == 4))? 1'd1 : 0;
  reg [32-1:0] _stream_avg_pool_serial_52_sink_5_sink_fsm_1;
  localparam _stream_avg_pool_serial_52_sink_5_sink_fsm_1_init = 0;
  wire _set_flag_1535;
  assign _set_flag_1535 = avg_pool_serial_52_comp_fsm == 5;
  assign _stream_avg_pool_serial_52_run_flag = (_set_flag_1535)? 1 : 0;
  reg _tmp_1536;
  reg _tmp_1537;
  reg _tmp_1538;
  reg _tmp_1539;
  reg _tmp_1540;
  reg _tmp_1541;
  reg _tmp_1542;
  reg _tmp_1543;
  reg _tmp_1544;
  reg _tmp_1545;
  assign _acc_0_source_stop = _acc_0_stream_oready && 1'd0;
  reg _tmp_1546;
  reg _tmp_1547;
  reg _tmp_1548;
  reg _tmp_1549;
  assign _acc_0_sink_start = _tmp_1549;
  reg _tmp_1550;
  reg _tmp_1551;
  reg _tmp_1552;
  reg _tmp_1553;
  assign _acc_0_sink_stop = _tmp_1553;
  reg _tmp_1554;
  reg _tmp_1555;
  reg _tmp_1556;
  reg _tmp_1557;
  assign _acc_0_sink_busy = _tmp_1557;
  reg _tmp_1558;
  assign _acc_0_busy = _acc_0_source_busy || _acc_0_sink_busy || _acc_0_busy_reg;
  reg _tmp_1559;
  reg _tmp_1560;
  reg _tmp_1561;
  reg _tmp_1562;
  reg _tmp_1563;
  reg _tmp_1564;
  reg [1-1:0] __variable_wdata_915;
  assign stream_avg_pool_serial_52__reduce_reset_data = __variable_wdata_915;
  reg _tmp_1565;
  reg _tmp_1566;
  reg _tmp_1567;
  reg _tmp_1568;
  assign _stream_avg_pool_serial_52_source_stop = _stream_avg_pool_serial_52_stream_oready && (_stream_avg_pool_serial_52_source_1_idle && (_stream_avg_pool_serial_52_fsm == 3));
  localparam _tmp_1569 = 1;
  wire [_tmp_1569-1:0] _tmp_1570;
  assign _tmp_1570 = _stream_avg_pool_serial_52_source_1_idle && (_stream_avg_pool_serial_52_fsm == 3);
  reg [_tmp_1569-1:0] _tmp_1571;
  localparam _tmp_1572 = 1;
  wire [_tmp_1572-1:0] _tmp_1573;
  assign _tmp_1573 = _stream_avg_pool_serial_52_source_1_idle && (_stream_avg_pool_serial_52_fsm == 3);
  reg [_tmp_1572-1:0] _tmp_1574;
  reg _tmp_1575;
  reg _tmp_1576;
  reg _tmp_1577;
  reg _tmp_1578;
  reg _tmp_1579;
  reg _tmp_1580;
  reg _tmp_1581;
  reg _tmp_1582;
  assign _stream_avg_pool_serial_52_sink_start = _tmp_1582;
  reg _tmp_1583;
  reg _tmp_1584;
  reg _tmp_1585;
  reg _tmp_1586;
  reg _tmp_1587;
  reg _tmp_1588;
  reg _tmp_1589;
  reg _tmp_1590;
  assign _stream_avg_pool_serial_52_sink_stop = _tmp_1590;
  reg _tmp_1591;
  reg _tmp_1592;
  reg _tmp_1593;
  reg _tmp_1594;
  reg _tmp_1595;
  reg _tmp_1596;
  reg _tmp_1597;
  reg _tmp_1598;
  assign _stream_avg_pool_serial_52_sink_busy = _tmp_1598;
  reg _tmp_1599;
  assign _stream_avg_pool_serial_52_busy = _stream_avg_pool_serial_52_source_busy || _stream_avg_pool_serial_52_sink_busy || _stream_avg_pool_serial_52_busy_reg;
  wire [12-1:0] _dma_write_packed_high_local_size_1600;
  assign _dma_write_packed_high_local_size_1600 = cparam_avg_pool_serial_52_out_write_size >> 2;
  wire [2-1:0] _dma_write_packed_low_local_size_1601;
  assign _dma_write_packed_low_local_size_1601 = cparam_avg_pool_serial_52_out_write_size & { 2{ 1'd1 } };
  wire [12-1:0] _dma_write_packed_local_packed_size_1602;
  assign _dma_write_packed_local_packed_size_1602 = (_dma_write_packed_low_local_size_1601 > 0)? _dma_write_packed_high_local_size_1600 + 1 : _dma_write_packed_high_local_size_1600;
  wire [32-1:0] mask_addr_shifted_1603;
  assign mask_addr_shifted_1603 = avg_pool_serial_52_objaddr + avg_pool_serial_52_out_base_offset + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_1604;
  assign mask_addr_masked_1604 = mask_addr_shifted_1603 << 2;
  reg [32-1:0] read_burst_packed_fsm_28;
  localparam read_burst_packed_fsm_28_init = 0;
  reg [14-1:0] read_burst_packed_addr_1605;
  reg [14-1:0] read_burst_packed_stride_1606;
  reg [33-1:0] read_burst_packed_length_1607;
  reg read_burst_packed_rvalid_1608;
  reg read_burst_packed_rlast_1609;
  wire [12-1:0] read_burst_packed_ram_addr_1610;
  assign read_burst_packed_ram_addr_1610 = read_burst_packed_addr_1605 >> 2;
  assign ram_w8_l16384_id1_0_1_addr = ((read_burst_packed_fsm_28 == 1) && (!read_burst_packed_rvalid_1608 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)))? read_burst_packed_ram_addr_1610 : 
                                      ((write_burst_packed_fsm_13 == 1) && write_burst_block_ram_wvalid_257)? write_burst_packed_ram_addr_263 : 'hx;
  assign ram_w8_l16384_id1_0_1_enable = ((read_burst_packed_fsm_28 == 1) && (!read_burst_packed_rvalid_1608 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)))? 1'd1 : 
                                        ((write_burst_packed_fsm_13 == 1) && write_burst_block_ram_wvalid_257)? 1'd1 : 0;
  localparam _tmp_1611 = 1;
  wire [_tmp_1611-1:0] _tmp_1612;
  assign _tmp_1612 = (read_burst_packed_fsm_28 == 1) && (!read_burst_packed_rvalid_1608 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0));
  reg [_tmp_1611-1:0] __tmp_1612_1;
  wire [8-1:0] read_burst_packed_ram_rdata_1613;
  assign read_burst_packed_ram_rdata_1613 = ram_w8_l16384_id1_0_1_rdata;
  wire [12-1:0] read_burst_packed_ram_addr_1614;
  assign read_burst_packed_ram_addr_1614 = read_burst_packed_addr_1605 >> 2;
  assign ram_w8_l16384_id1_1_1_addr = ((read_burst_packed_fsm_28 == 1) && (!read_burst_packed_rvalid_1608 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)))? read_burst_packed_ram_addr_1614 : 
                                      ((write_burst_packed_fsm_13 == 1) && write_burst_block_ram_wvalid_257)? write_burst_packed_ram_addr_265 : 'hx;
  assign ram_w8_l16384_id1_1_1_enable = ((read_burst_packed_fsm_28 == 1) && (!read_burst_packed_rvalid_1608 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)))? 1'd1 : 
                                        ((write_burst_packed_fsm_13 == 1) && write_burst_block_ram_wvalid_257)? 1'd1 : 0;
  localparam _tmp_1615 = 1;
  wire [_tmp_1615-1:0] _tmp_1616;
  assign _tmp_1616 = (read_burst_packed_fsm_28 == 1) && (!read_burst_packed_rvalid_1608 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0));
  reg [_tmp_1615-1:0] __tmp_1616_1;
  wire [8-1:0] read_burst_packed_ram_rdata_1617;
  assign read_burst_packed_ram_rdata_1617 = ram_w8_l16384_id1_1_1_rdata;
  wire [12-1:0] read_burst_packed_ram_addr_1618;
  assign read_burst_packed_ram_addr_1618 = read_burst_packed_addr_1605 >> 2;
  assign ram_w8_l16384_id1_2_1_addr = ((read_burst_packed_fsm_28 == 1) && (!read_burst_packed_rvalid_1608 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)))? read_burst_packed_ram_addr_1618 : 
                                      ((write_burst_packed_fsm_13 == 1) && write_burst_block_ram_wvalid_257)? write_burst_packed_ram_addr_267 : 'hx;
  assign ram_w8_l16384_id1_2_1_enable = ((read_burst_packed_fsm_28 == 1) && (!read_burst_packed_rvalid_1608 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)))? 1'd1 : 
                                        ((write_burst_packed_fsm_13 == 1) && write_burst_block_ram_wvalid_257)? 1'd1 : 0;
  localparam _tmp_1619 = 1;
  wire [_tmp_1619-1:0] _tmp_1620;
  assign _tmp_1620 = (read_burst_packed_fsm_28 == 1) && (!read_burst_packed_rvalid_1608 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0));
  reg [_tmp_1619-1:0] __tmp_1620_1;
  wire [8-1:0] read_burst_packed_ram_rdata_1621;
  assign read_burst_packed_ram_rdata_1621 = ram_w8_l16384_id1_2_1_rdata;
  wire [12-1:0] read_burst_packed_ram_addr_1622;
  assign read_burst_packed_ram_addr_1622 = read_burst_packed_addr_1605 >> 2;
  assign ram_w8_l16384_id1_3_1_addr = ((read_burst_packed_fsm_28 == 1) && (!read_burst_packed_rvalid_1608 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)))? read_burst_packed_ram_addr_1622 : 
                                      ((write_burst_packed_fsm_13 == 1) && write_burst_block_ram_wvalid_257)? write_burst_packed_ram_addr_269 : 'hx;
  assign ram_w8_l16384_id1_3_1_enable = ((read_burst_packed_fsm_28 == 1) && (!read_burst_packed_rvalid_1608 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)))? 1'd1 : 
                                        ((write_burst_packed_fsm_13 == 1) && write_burst_block_ram_wvalid_257)? 1'd1 : 0;
  localparam _tmp_1623 = 1;
  wire [_tmp_1623-1:0] _tmp_1624;
  assign _tmp_1624 = (read_burst_packed_fsm_28 == 1) && (!read_burst_packed_rvalid_1608 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0));
  reg [_tmp_1623-1:0] __tmp_1624_1;
  wire [8-1:0] read_burst_packed_ram_rdata_1625;
  assign read_burst_packed_ram_rdata_1625 = ram_w8_l16384_id1_3_1_rdata;
  wire [32-1:0] read_burst_packed_rdata_1626;
  assign read_burst_packed_rdata_1626 = { read_burst_packed_ram_rdata_1625, read_burst_packed_ram_rdata_1621, read_burst_packed_ram_rdata_1617, read_burst_packed_ram_rdata_1613 };
  assign _maxi_write_req_fifo_deq = ((_maxi_write_data_fsm == 2) && (!_maxi_write_req_fifo_empty && (_maxi_write_size_buf == 0)) && !_maxi_write_req_fifo_empty)? 1 : 
                                    ((_maxi_write_data_fsm == 0) && (!_maxi_write_data_busy && !_maxi_write_req_fifo_empty && (_maxi_write_op_sel_fifo == 3)) && !_maxi_write_req_fifo_empty)? 1 : 
                                    ((_maxi_write_data_fsm == 2) && (!_maxi_write_req_fifo_empty && (_maxi_write_size_buf == 0)) && !_maxi_write_req_fifo_empty)? 1 : 
                                    ((_maxi_write_data_fsm == 0) && (!_maxi_write_data_busy && !_maxi_write_req_fifo_empty && (_maxi_write_op_sel_fifo == 2)) && !_maxi_write_req_fifo_empty)? 1 : 
                                    ((_maxi_write_data_fsm == 2) && (!_maxi_write_req_fifo_empty && (_maxi_write_size_buf == 0)) && !_maxi_write_req_fifo_empty)? 1 : 
                                    ((_maxi_write_data_fsm == 0) && (!_maxi_write_data_busy && !_maxi_write_req_fifo_empty && (_maxi_write_op_sel_fifo == 1)) && !_maxi_write_req_fifo_empty)? 1 : 0;
  reg _maxi_wdata_cond_2_1;
  reg [32-1:0] matmul_55_objaddr;
  reg [32-1:0] matmul_55_arg_objaddr_0;
  reg [32-1:0] matmul_55_arg_objaddr_1;
  reg [32-1:0] matmul_55_arg_objaddr_2;
  reg [32-1:0] matmul_55_arg_objaddr_3;
  reg [32-1:0] control_matmul_55;
  localparam control_matmul_55_init = 0;
  reg _control_matmul_55_called;
  wire signed [32-1:0] matmul_55_act_base_offset;
  reg signed [32-1:0] matmul_55_act_base_offset_row;
  reg signed [32-1:0] matmul_55_act_base_offset_bat;
  assign matmul_55_act_base_offset = matmul_55_act_base_offset_row + matmul_55_act_base_offset_bat;
  reg signed [32-1:0] matmul_55_filter_base_offset;
  reg [32-1:0] matmul_55_next_stream_num_ops;
  wire signed [32-1:0] matmul_55_out_base_offset;
  reg signed [32-1:0] matmul_55_out_base_offset_val;
  reg signed [32-1:0] matmul_55_out_base_offset_col;
  reg signed [32-1:0] matmul_55_out_base_offset_row;
  reg signed [32-1:0] matmul_55_out_base_offset_bat;
  reg signed [32-1:0] matmul_55_out_base_offset_och;
  assign matmul_55_out_base_offset = matmul_55_out_base_offset_val + matmul_55_out_base_offset_col + matmul_55_out_base_offset_row + matmul_55_out_base_offset_bat + matmul_55_out_base_offset_och;
  reg matmul_55_dma_flag_0;
  reg [32-1:0] matmul_55_sync_comp_count;
  reg [32-1:0] matmul_55_sync_out_count;
  reg [32-1:0] matmul_55_write_count;
  reg [32-1:0] matmul_55_next_out_write_size;
  reg [32-1:0] matmul_55_col_count;
  reg [32-1:0] matmul_55_row_count;
  reg [32-1:0] matmul_55_bat_count;
  reg [32-1:0] matmul_55_och_count;
  reg [1-1:0] matmul_55_col_select;
  reg [1-1:0] matmul_55_row_select;
  reg [32-1:0] matmul_55_out_col_count;
  reg [32-1:0] matmul_55_out_row_count;
  reg [32-1:0] matmul_55_out_ram_select;
  reg [32-1:0] matmul_55_prev_col_count;
  reg [32-1:0] matmul_55_prev_row_count;
  reg [32-1:0] matmul_55_prev_bat_count;
  reg [32-1:0] matmul_55_prev_och_count;
  reg [1-1:0] matmul_55_prev_row_select;
  reg [32-1:0] matmul_55_stream_act_local_0;
  reg [32-1:0] matmul_55_stream_out_local_val;
  reg [32-1:0] matmul_55_stream_out_local_col;
  wire [32-1:0] matmul_55_stream_out_local;
  assign matmul_55_stream_out_local = matmul_55_stream_out_local_val + matmul_55_stream_out_local_col;
  reg [32-1:0] matmul_55_act_page_comp_offset_0;
  reg [32-1:0] matmul_55_act_page_dma_offset_0;
  reg [32-1:0] matmul_55_filter_page_comp_offset;
  reg [32-1:0] matmul_55_filter_page_dma_offset;
  reg matmul_55_out_page;
  reg [32-1:0] matmul_55_out_page_comp_offset;
  reg [32-1:0] matmul_55_out_page_dma_offset;
  reg [32-1:0] matmul_55_out_laddr_offset;
  reg matmul_55_skip_read_filter;
  reg matmul_55_skip_read_act;
  reg matmul_55_skip_comp;
  reg matmul_55_skip_write_out;
  wire [32-1:0] mask_addr_shifted_1627;
  assign mask_addr_shifted_1627 = matmul_55_arg_objaddr_2 + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_1628;
  assign mask_addr_masked_1628 = mask_addr_shifted_1627 << 2;
  wire [1-1:0] _dma_read_packed_high_local_size_1629;
  assign _dma_read_packed_high_local_size_1629 = cparam_matmul_55_scale_num >> 2;
  wire [2-1:0] _dma_read_packed_low_local_size_1630;
  assign _dma_read_packed_low_local_size_1630 = cparam_matmul_55_scale_num & { 2{ 1'd1 } };
  wire [1-1:0] _dma_read_packed_local_packed_size_1631;
  assign _dma_read_packed_local_packed_size_1631 = (_dma_read_packed_low_local_size_1630 > 0)? _dma_read_packed_high_local_size_1629 + 1 : _dma_read_packed_high_local_size_1629;
  wire [32-1:0] mask_addr_shifted_1632;
  assign mask_addr_shifted_1632 = matmul_55_arg_objaddr_3 + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_1633;
  assign mask_addr_masked_1633 = mask_addr_shifted_1632 << 2;
  wire [18-1:0] _dma_read_packed_high_local_size_1634;
  assign _dma_read_packed_high_local_size_1634 = cparam_matmul_55_filter_read_size >> 2;
  wire [2-1:0] _dma_read_packed_low_local_size_1635;
  assign _dma_read_packed_low_local_size_1635 = cparam_matmul_55_filter_read_size & { 2{ 1'd1 } };
  wire [18-1:0] _dma_read_packed_local_packed_size_1636;
  assign _dma_read_packed_local_packed_size_1636 = (_dma_read_packed_low_local_size_1635 > 0)? _dma_read_packed_high_local_size_1634 + 1 : _dma_read_packed_high_local_size_1634;
  wire [32-1:0] mask_addr_shifted_1637;
  assign mask_addr_shifted_1637 = matmul_55_arg_objaddr_1 + matmul_55_filter_base_offset + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_1638;
  assign mask_addr_masked_1638 = mask_addr_shifted_1637 << 2;
  wire [32-1:0] matmul_55_mux_act_gaddr_0;
  assign matmul_55_mux_act_gaddr_0 = (matmul_55_row_select == 0)? matmul_55_arg_objaddr_0 + (matmul_55_act_base_offset + cparam_matmul_55_act_offset_values_0) : 1'd0;
  wire matmul_55_dma_pad_mask_0;
  assign matmul_55_dma_pad_mask_0 = (matmul_55_row_count + 0 < cparam_matmul_55_pad_row_top) || (matmul_55_row_count + 0 >= cparam_matmul_55_act_num_row + cparam_matmul_55_pad_row_top);
  wire matmul_55_mux_dma_pad_mask_0;
  assign matmul_55_mux_dma_pad_mask_0 = (matmul_55_row_select == 0)? matmul_55_dma_pad_mask_0 : 1'd0;
  wire matmul_55_mux_dma_flag_0;
  assign matmul_55_mux_dma_flag_0 = (matmul_55_prev_row_select == 0)? matmul_55_dma_flag_0 : 1'd0;
  wire [15-1:0] _dma_read_packed_high_local_size_1639;
  assign _dma_read_packed_high_local_size_1639 = cparam_matmul_55_act_read_size >> 2;
  wire [2-1:0] _dma_read_packed_low_local_size_1640;
  assign _dma_read_packed_low_local_size_1640 = cparam_matmul_55_act_read_size & { 2{ 1'd1 } };
  wire [15-1:0] _dma_read_packed_local_packed_size_1641;
  assign _dma_read_packed_local_packed_size_1641 = (_dma_read_packed_low_local_size_1640 > 0)? _dma_read_packed_high_local_size_1639 + 1 : _dma_read_packed_high_local_size_1639;
  wire [32-1:0] mask_addr_shifted_1642;
  assign mask_addr_shifted_1642 = matmul_55_mux_act_gaddr_0 + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_1643;
  assign mask_addr_masked_1643 = mask_addr_shifted_1642 << 2;
  assign _maxi_read_req_fifo_deq = ((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 9)) && !_maxi_read_req_fifo_empty)? 1 : 
                                   ((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 8)) && !_maxi_read_req_fifo_empty)? 1 : 
                                   ((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 7)) && !_maxi_read_req_fifo_empty)? 1 : 
                                   ((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 6)) && !_maxi_read_req_fifo_empty)? 1 : 
                                   ((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 5)) && !_maxi_read_req_fifo_empty)? 1 : 
                                   ((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 4)) && !_maxi_read_req_fifo_empty)? 1 : 
                                   ((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 3)) && !_maxi_read_req_fifo_empty)? 1 : 
                                   ((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 2)) && !_maxi_read_req_fifo_empty)? 1 : 
                                   ((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 1)) && !_maxi_read_req_fifo_empty)? 1 : 0;
  reg [32-1:0] write_burst_packed_fsm_29;
  localparam write_burst_packed_fsm_29_init = 0;
  reg [15-1:0] write_burst_packed_addr_1644;
  reg [15-1:0] write_burst_packed_stride_1645;
  reg [33-1:0] write_burst_packed_length_1646;
  reg write_burst_packed_done_1647;
  wire [13-1:0] write_burst_packed_ram_addr_1648;
  assign write_burst_packed_ram_addr_1648 = write_burst_packed_addr_1644 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_1649;
  assign write_burst_packed_ram_wdata_1649 = _maxi_rdata_sb_0 >> 0;
  assign ram_w8_l32768_id0_0_1_addr = ((write_burst_packed_fsm_29 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_addr_1648 : 'hx;
  assign ram_w8_l32768_id0_0_1_wdata = ((write_burst_packed_fsm_29 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_wdata_1649 : 'hx;
  assign ram_w8_l32768_id0_0_1_wenable = ((write_burst_packed_fsm_29 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  assign ram_w8_l32768_id0_0_1_enable = ((write_burst_packed_fsm_29 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  wire [13-1:0] write_burst_packed_ram_addr_1650;
  assign write_burst_packed_ram_addr_1650 = write_burst_packed_addr_1644 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_1651;
  assign write_burst_packed_ram_wdata_1651 = _maxi_rdata_sb_0 >> 8;
  assign ram_w8_l32768_id0_1_1_addr = ((write_burst_packed_fsm_29 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_addr_1650 : 'hx;
  assign ram_w8_l32768_id0_1_1_wdata = ((write_burst_packed_fsm_29 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_wdata_1651 : 'hx;
  assign ram_w8_l32768_id0_1_1_wenable = ((write_burst_packed_fsm_29 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  assign ram_w8_l32768_id0_1_1_enable = ((write_burst_packed_fsm_29 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  wire [13-1:0] write_burst_packed_ram_addr_1652;
  assign write_burst_packed_ram_addr_1652 = write_burst_packed_addr_1644 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_1653;
  assign write_burst_packed_ram_wdata_1653 = _maxi_rdata_sb_0 >> 16;
  assign ram_w8_l32768_id0_2_1_addr = ((write_burst_packed_fsm_29 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_addr_1652 : 'hx;
  assign ram_w8_l32768_id0_2_1_wdata = ((write_burst_packed_fsm_29 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_wdata_1653 : 'hx;
  assign ram_w8_l32768_id0_2_1_wenable = ((write_burst_packed_fsm_29 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  assign ram_w8_l32768_id0_2_1_enable = ((write_burst_packed_fsm_29 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  wire [13-1:0] write_burst_packed_ram_addr_1654;
  assign write_burst_packed_ram_addr_1654 = write_burst_packed_addr_1644 >> 2;
  wire [8-1:0] write_burst_packed_ram_wdata_1655;
  assign write_burst_packed_ram_wdata_1655 = _maxi_rdata_sb_0 >> 24;
  assign ram_w8_l32768_id0_3_1_addr = ((write_burst_packed_fsm_29 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_addr_1654 : 'hx;
  assign ram_w8_l32768_id0_3_1_wdata = ((write_burst_packed_fsm_29 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_wdata_1655 : 'hx;
  assign ram_w8_l32768_id0_3_1_wenable = ((write_burst_packed_fsm_29 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  assign ram_w8_l32768_id0_3_1_enable = ((write_burst_packed_fsm_29 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  assign _maxi_rready_sb_0 = (_maxi_read_data_fsm == 2) || (_maxi_read_data_fsm == 2) || (_maxi_read_data_fsm == 2) || (_maxi_read_data_fsm == 2) || (_maxi_read_data_fsm == 2) || (_maxi_read_data_fsm == 2) || (_maxi_read_data_fsm == 2) || (_maxi_read_data_fsm == 2) || (_maxi_read_data_fsm == 2);
  reg [32-1:0] matmul_55_comp_fsm;
  localparam matmul_55_comp_fsm_init = 0;
  reg [32-1:0] matmul_55_filter_page_comp_offset_buf;
  reg [32-1:0] matmul_55_act_page_comp_offset_buf_0;
  reg [32-1:0] matmul_55_out_page_comp_offset_buf;
  reg [32-1:0] matmul_55_row_count_buf;
  reg [1-1:0] matmul_55_row_select_buf;
  reg [32-1:0] matmul_55_och_count_buf;
  wire matmul_55_stream_pad_mask_0_0;
  assign matmul_55_stream_pad_mask_0_0 = (matmul_55_col_count + 0 < cparam_matmul_55_pad_col_left) || (matmul_55_col_count + 0 >= cparam_matmul_55_act_num_col + cparam_matmul_55_pad_col_left) || (matmul_55_row_count_buf + 0 < cparam_matmul_55_pad_row_top) || (matmul_55_row_count_buf + 0 >= cparam_matmul_55_act_num_row + cparam_matmul_55_pad_row_top);
  reg [1-1:0] matmul_55_stream_pad_masks;
  wire [15-1:0] stream_matmul_55_parameter_0_data;
  wire [1-1:0] stream_matmul_55_parameter_1_data;
  wire [1-1:0] stream_matmul_55_parameter_2_data;
  wire [1-1:0] stream_matmul_55_parameter_3_data;
  wire [1-1:0] stream_matmul_55_parameter_4_data;
  wire [1-1:0] stream_matmul_55__reduce_reset_data;
  wire [1-1:0] stream_matmul_55_parameter_6_data;
  wire [32-1:0] stream_matmul_55_source_7_data;
  wire [1-1:0] stream_matmul_55_parameter_8_data;
  wire [8-1:0] stream_matmul_55_source_9_data;
  wire [1-1:0] stream_matmul_55_parameter_10_data;
  wire [8-1:0] stream_matmul_55_source_11_data;
  wire [1-1:0] stream_matmul_55_parameter_12_data;
  wire [8-1:0] stream_matmul_55_source_13_data;
  wire [1-1:0] stream_matmul_55_parameter_14_data;
  wire [8-1:0] stream_matmul_55_source_15_data;
  wire [1-1:0] stream_matmul_55_parameter_16_data;
  wire [1-1:0] stream_matmul_55_parameter_17_data;
  wire [5-1:0] stream_matmul_55_parameter_18_data;
  wire [2-1:0] stream_matmul_55_parameter_19_data;
  wire [8-1:0] stream_matmul_55_source_20_data;
  wire [8-1:0] stream_matmul_55_source_21_data;
  reg __stream_matmul_55_stream_ivalid_1;
  reg __stream_matmul_55_stream_ivalid_2;
  reg __stream_matmul_55_stream_ivalid_3;
  reg __stream_matmul_55_stream_ivalid_4;
  reg __stream_matmul_55_stream_ivalid_5;
  reg __stream_matmul_55_stream_ivalid_6;
  reg __stream_matmul_55_stream_ivalid_7;
  reg __stream_matmul_55_stream_ivalid_8;
  reg __stream_matmul_55_stream_ivalid_9;
  reg __stream_matmul_55_stream_ivalid_10;
  reg __stream_matmul_55_stream_ivalid_11;
  reg __stream_matmul_55_stream_ivalid_12;
  reg __stream_matmul_55_stream_ivalid_13;
  reg __stream_matmul_55_stream_ivalid_14;
  reg __stream_matmul_55_stream_ivalid_15;
  reg __stream_matmul_55_stream_ivalid_16;
  reg __stream_matmul_55_stream_ivalid_17;
  reg __stream_matmul_55_stream_ivalid_18;
  reg __stream_matmul_55_stream_ivalid_19;
  reg __stream_matmul_55_stream_ivalid_20;
  reg __stream_matmul_55_stream_ivalid_21;
  reg __stream_matmul_55_stream_ivalid_22;
  reg __stream_matmul_55_stream_ivalid_23;
  reg __stream_matmul_55_stream_ivalid_24;
  reg __stream_matmul_55_stream_ivalid_25;
  reg __stream_matmul_55_stream_ivalid_26;
  reg __stream_matmul_55_stream_ivalid_27;
  reg __stream_matmul_55_stream_ivalid_28;
  reg __stream_matmul_55_stream_ivalid_29;
  wire [32-1:0] _slice_data_955;
  assign _slice_data_955 = stream_matmul_55_source_7_data[6'd31:1'd0];
  wire [32-1:0] _reinterpretcast_src_956;
  assign _reinterpretcast_src_956 = _slice_data_955;
  wire signed [32-1:0] _reinterpretcast_data_956;
  assign _reinterpretcast_data_956 = _reinterpretcast_src_956;
  wire signed [32-1:0] _cond_data_957;
  assign _cond_data_957 = (stream_matmul_55_parameter_6_data)? _reinterpretcast_data_956 : _reinterpretcast_data_956;
  wire [8-1:0] _slice_data_962;
  assign _slice_data_962 = stream_matmul_55_source_9_data[4'd7:1'd0];
  wire [8-1:0] _reinterpretcast_src_963;
  assign _reinterpretcast_src_963 = _slice_data_962;
  wire signed [8-1:0] _reinterpretcast_data_963;
  assign _reinterpretcast_data_963 = _reinterpretcast_src_963;
  wire signed [8-1:0] _cond_data_964;
  assign _cond_data_964 = (stream_matmul_55_parameter_8_data)? _reinterpretcast_data_963 : _reinterpretcast_data_963;
  wire [8-1:0] _slice_data_969;
  assign _slice_data_969 = stream_matmul_55_source_11_data[4'd7:1'd0];
  wire [8-1:0] _reinterpretcast_src_970;
  assign _reinterpretcast_src_970 = _slice_data_969;
  wire [8-1:0] _reinterpretcast_data_970;
  assign _reinterpretcast_data_970 = _reinterpretcast_src_970;
  wire [8-1:0] _cond_data_971;
  assign _cond_data_971 = (stream_matmul_55_parameter_10_data)? _reinterpretcast_data_970 : _reinterpretcast_data_970;
  wire [8-1:0] _slice_data_976;
  assign _slice_data_976 = stream_matmul_55_source_13_data[4'd7:1'd0];
  wire [8-1:0] _reinterpretcast_src_977;
  assign _reinterpretcast_src_977 = _slice_data_976;
  wire [8-1:0] _reinterpretcast_data_977;
  assign _reinterpretcast_data_977 = _reinterpretcast_src_977;
  wire [8-1:0] _cond_data_978;
  assign _cond_data_978 = (stream_matmul_55_parameter_12_data)? _reinterpretcast_data_977 : _reinterpretcast_data_977;
  wire [8-1:0] _slice_data_983;
  assign _slice_data_983 = stream_matmul_55_source_15_data[4'd7:1'd0];
  wire [8-1:0] _reinterpretcast_src_984;
  assign _reinterpretcast_src_984 = _slice_data_983;
  wire [8-1:0] _reinterpretcast_data_984;
  assign _reinterpretcast_data_984 = _reinterpretcast_src_984;
  wire [8-1:0] _cond_data_985;
  assign _cond_data_985 = (stream_matmul_55_parameter_14_data)? _reinterpretcast_data_984 : _reinterpretcast_data_984;
  reg [1-1:0] _eq_data_991;
  reg [1-1:0] _eq_data_995;
  wire [8-1:0] _reinterpretcast_src_1009;
  assign _reinterpretcast_src_1009 = stream_matmul_55_source_21_data;
  wire signed [8-1:0] _reinterpretcast_data_1009;
  assign _reinterpretcast_data_1009 = _reinterpretcast_src_1009;
  wire [1-1:0] _pointer_data_1010;
  assign _pointer_data_1010 = stream_matmul_55_parameter_3_data[1'sd0];
  reg [8-1:0] _plus_data_1015;
  reg [8-1:0] _plus_data_1020;
  reg [8-1:0] _plus_data_1025;
  reg [1-1:0] _eq_data_1031;
  reg [1-1:0] _eq_data_1034;
  reg [8-1:0] __delay_data_1192__variable_990;
  reg [1-1:0] __delay_data_1193_pointer_1010;
  reg signed [8-1:0] __delay_data_1194_reinterpretcast_1009;
  reg [1-1:0] __delay_data_1195__variable_941;
  reg [15-1:0] __delay_data_1216__variable_936;
  reg signed [32-1:0] __delay_data_1227_cond_957;
  reg signed [8-1:0] __delay_data_1244_cond_964;
  wire signed [8-1:0] _cond_data_993;
  assign _cond_data_993 = (_eq_data_991)? __delay_data_1192__variable_990 : 1'sd0;
  wire signed [8-1:0] _cond_data_997;
  assign _cond_data_997 = (_eq_data_995)? _cond_data_993 : 1'sd0;
  wire signed [8-1:0] _reinterpretcast_src_1003;
  assign _reinterpretcast_src_1003 = _cond_data_997;
  wire signed [8-1:0] _reinterpretcast_data_1003;
  assign _reinterpretcast_data_1003 = _reinterpretcast_src_1003;
  wire signed [8-1:0] _cond_data_1013;
  assign _cond_data_1013 = (__delay_data_1193_pointer_1010)? 1'sd0 : _reinterpretcast_data_1003;
  assign _mul_5_is_root = ((_stream_matmul_55_busy)? 0 : 1) && (((_stream_conv2d_24_busy)? 0 : 1) && 1);
  assign _mul_5_stream_oready = ((_stream_matmul_55_busy)? _stream_matmul_55_stream_oready : 1) && (((_stream_conv2d_24_busy)? _stream_conv2d_24_stream_oready : 1) && _mul_5_stream_internal_oready);
  reg [1-1:0] __delay_data_1196__delay_1195__variable_941;
  reg [8-1:0] __delay_data_1206_plus_1020;
  reg [15-1:0] __delay_data_1217__delay_1216__variable_936;
  reg signed [32-1:0] __delay_data_1228__delay_1227_cond_957;
  reg signed [8-1:0] __delay_data_1245__delay_1244_cond_964;
  reg [8-1:0] __delay_data_1262_plus_1025;
  reg [1-1:0] __delay_data_1280_eq_1031;
  reg [1-1:0] __delay_data_1309_eq_1034;
  reg [1-1:0] __delay_data_1197__delay_1196__delay_1195__variable_941;
  reg [8-1:0] __delay_data_1207__delay_1206_plus_1020;
  reg [15-1:0] __delay_data_1218__delay_1217__delay_1216__variable_936;
  reg signed [32-1:0] __delay_data_1229__delay_1228__delay_1227_cond_957;
  reg signed [8-1:0] __delay_data_1246__delay_1245__delay_1244_cond_964;
  reg [8-1:0] __delay_data_1263__delay_1262_plus_1025;
  reg [1-1:0] __delay_data_1281__delay_1280_eq_1031;
  reg [1-1:0] __delay_data_1310__delay_1309_eq_1034;
  reg [1-1:0] __delay_data_1198__delay_1197__delay_1196____variable_941;
  reg [8-1:0] __delay_data_1208__delay_1207__delay_1206_plus_1020;
  reg [15-1:0] __delay_data_1219__delay_1218__delay_1217____variable_936;
  reg signed [32-1:0] __delay_data_1230__delay_1229__delay_1228__delay_1227_cond_957;
  reg signed [8-1:0] __delay_data_1247__delay_1246__delay_1245__delay_1244_cond_964;
  reg [8-1:0] __delay_data_1264__delay_1263__delay_1262_plus_1025;
  reg [1-1:0] __delay_data_1282__delay_1281__delay_1280_eq_1031;
  reg [1-1:0] __delay_data_1311__delay_1310__delay_1309_eq_1034;
  reg [1-1:0] __delay_data_1199__delay_1198__delay_1197____variable_941;
  reg [8-1:0] __delay_data_1209__delay_1208__delay_1207___plus_1020;
  reg [15-1:0] __delay_data_1220__delay_1219__delay_1218____variable_936;
  reg signed [32-1:0] __delay_data_1231__delay_1230__delay_1229__delay_1228___cond_957;
  reg signed [8-1:0] __delay_data_1248__delay_1247__delay_1246__delay_1245___cond_964;
  reg [8-1:0] __delay_data_1265__delay_1264__delay_1263___plus_1025;
  reg [1-1:0] __delay_data_1283__delay_1282__delay_1281__delay_1280_eq_1031;
  reg [1-1:0] __delay_data_1312__delay_1311__delay_1310__delay_1309_eq_1034;
  reg [1-1:0] __delay_data_1200__delay_1199__delay_1198____variable_941;
  reg [8-1:0] __delay_data_1210__delay_1209__delay_1208___plus_1020;
  reg [15-1:0] __delay_data_1221__delay_1220__delay_1219____variable_936;
  reg signed [32-1:0] __delay_data_1232__delay_1231__delay_1230__delay_1229___cond_957;
  reg signed [8-1:0] __delay_data_1249__delay_1248__delay_1247__delay_1246___cond_964;
  reg [8-1:0] __delay_data_1266__delay_1265__delay_1264___plus_1025;
  reg [1-1:0] __delay_data_1284__delay_1283__delay_1282__delay_1281___eq_1031;
  reg [1-1:0] __delay_data_1313__delay_1312__delay_1311__delay_1310___eq_1034;
  reg [1-1:0] __delay_data_1201__delay_1200__delay_1199____variable_941;
  reg [8-1:0] __delay_data_1211__delay_1210__delay_1209___plus_1020;
  reg [15-1:0] __delay_data_1222__delay_1221__delay_1220____variable_936;
  reg signed [32-1:0] __delay_data_1233__delay_1232__delay_1231__delay_1230___cond_957;
  reg signed [8-1:0] __delay_data_1250__delay_1249__delay_1248__delay_1247___cond_964;
  reg [8-1:0] __delay_data_1267__delay_1266__delay_1265___plus_1025;
  reg [1-1:0] __delay_data_1285__delay_1284__delay_1283__delay_1282___eq_1031;
  reg [1-1:0] __delay_data_1314__delay_1313__delay_1312__delay_1311___eq_1034;
  reg [1-1:0] __delay_data_1202__delay_1201__delay_1200____variable_941;
  reg [8-1:0] __delay_data_1212__delay_1211__delay_1210___plus_1020;
  reg [15-1:0] __delay_data_1223__delay_1222__delay_1221____variable_936;
  reg signed [32-1:0] __delay_data_1234__delay_1233__delay_1232__delay_1231___cond_957;
  reg signed [8-1:0] __delay_data_1251__delay_1250__delay_1249__delay_1248___cond_964;
  reg [8-1:0] __delay_data_1268__delay_1267__delay_1266___plus_1025;
  reg [1-1:0] __delay_data_1286__delay_1285__delay_1284__delay_1283___eq_1031;
  reg [1-1:0] __delay_data_1315__delay_1314__delay_1313__delay_1312___eq_1034;
  reg [1-1:0] __delay_data_1203__delay_1202__delay_1201____variable_941;
  reg [8-1:0] __delay_data_1213__delay_1212__delay_1211___plus_1020;
  reg [15-1:0] __delay_data_1224__delay_1223__delay_1222____variable_936;
  reg signed [32-1:0] __delay_data_1235__delay_1234__delay_1233__delay_1232___cond_957;
  reg signed [8-1:0] __delay_data_1252__delay_1251__delay_1250__delay_1249___cond_964;
  reg [8-1:0] __delay_data_1269__delay_1268__delay_1267___plus_1025;
  reg [1-1:0] __delay_data_1287__delay_1286__delay_1285__delay_1284___eq_1031;
  reg [1-1:0] __delay_data_1316__delay_1315__delay_1314__delay_1313___eq_1034;
  reg [1-1:0] __delay_data_1204__delay_1203__delay_1202____variable_941;
  reg [8-1:0] __delay_data_1214__delay_1213__delay_1212___plus_1020;
  reg [15-1:0] __delay_data_1225__delay_1224__delay_1223____variable_936;
  reg signed [32-1:0] __delay_data_1236__delay_1235__delay_1234__delay_1233___cond_957;
  reg signed [8-1:0] __delay_data_1253__delay_1252__delay_1251__delay_1250___cond_964;
  reg [8-1:0] __delay_data_1270__delay_1269__delay_1268___plus_1025;
  reg [1-1:0] __delay_data_1288__delay_1287__delay_1286__delay_1285___eq_1031;
  reg [1-1:0] __delay_data_1317__delay_1316__delay_1315__delay_1314___eq_1034;
  wire signed [16-1:0] __substreamoutput_data_1016;
  assign __substreamoutput_data_1016 = mul_5_z_data;
  reg signed [32-1:0] __variable_wdata_58;
  assign add_tree_2_var0_data = __variable_wdata_58;
  assign _add_tree_2_is_root = ((_stream_matmul_55_busy)? 0 : 1) && 1;
  assign _add_tree_2_stream_oready = ((_stream_matmul_55_busy)? _stream_matmul_55_stream_oready : 1) && _add_tree_2_stream_internal_oready;
  reg [1-1:0] __delay_data_1205__delay_1204__delay_1203____variable_941;
  reg [8-1:0] __delay_data_1215__delay_1214__delay_1213___plus_1020;
  reg [15-1:0] __delay_data_1226__delay_1225__delay_1224____variable_936;
  reg signed [32-1:0] __delay_data_1237__delay_1236__delay_1235__delay_1234___cond_957;
  reg signed [8-1:0] __delay_data_1254__delay_1253__delay_1252__delay_1251___cond_964;
  reg [8-1:0] __delay_data_1271__delay_1270__delay_1269___plus_1025;
  reg [1-1:0] __delay_data_1289__delay_1288__delay_1287__delay_1286___eq_1031;
  reg [1-1:0] __delay_data_1318__delay_1317__delay_1316__delay_1315___eq_1034;
  wire signed [32-1:0] __substreamoutput_data_1018;
  assign __substreamoutput_data_1018 = add_tree_2_sum_data;
  assign _acc_1_is_root = ((_stream_matmul_55_busy)? 0 : 1) && (((_stream_conv2d_24_busy)? 0 : 1) && 1);
  assign _acc_1_stream_oready = ((_stream_matmul_55_busy)? _stream_matmul_55_stream_oready : 1) && (((_stream_conv2d_24_busy)? _stream_conv2d_24_stream_oready : 1) && _acc_1_stream_internal_oready);
  reg signed [32-1:0] __delay_data_1238__delay_1237__delay_1236__delay_1235___cond_957;
  reg signed [8-1:0] __delay_data_1255__delay_1254__delay_1253__delay_1252___cond_964;
  reg [8-1:0] __delay_data_1272__delay_1271__delay_1270___plus_1025;
  reg [1-1:0] __delay_data_1290__delay_1289__delay_1288__delay_1287___eq_1031;
  reg [1-1:0] __delay_data_1319__delay_1318__delay_1317__delay_1316___eq_1034;
  reg signed [32-1:0] __delay_data_1239__delay_1238__delay_1237__delay_1236___cond_957;
  reg signed [8-1:0] __delay_data_1256__delay_1255__delay_1254__delay_1253___cond_964;
  reg [8-1:0] __delay_data_1273__delay_1272__delay_1271___plus_1025;
  reg [1-1:0] __delay_data_1291__delay_1290__delay_1289__delay_1288___eq_1031;
  reg [1-1:0] __delay_data_1320__delay_1319__delay_1318__delay_1317___eq_1034;
  reg signed [32-1:0] __delay_data_1240__delay_1239__delay_1238__delay_1237___cond_957;
  reg signed [8-1:0] __delay_data_1257__delay_1256__delay_1255__delay_1254___cond_964;
  reg [8-1:0] __delay_data_1274__delay_1273__delay_1272___plus_1025;
  reg [1-1:0] __delay_data_1292__delay_1291__delay_1290__delay_1289___eq_1031;
  reg [1-1:0] __delay_data_1321__delay_1320__delay_1319__delay_1318___eq_1034;
  reg signed [32-1:0] __delay_data_1241__delay_1240__delay_1239__delay_1238___cond_957;
  reg signed [8-1:0] __delay_data_1258__delay_1257__delay_1256__delay_1255___cond_964;
  reg [8-1:0] __delay_data_1275__delay_1274__delay_1273___plus_1025;
  reg [1-1:0] __delay_data_1293__delay_1292__delay_1291__delay_1290___eq_1031;
  reg [1-1:0] __delay_data_1322__delay_1321__delay_1320__delay_1319___eq_1034;
  reg signed [32-1:0] __delay_data_1242__delay_1241__delay_1240__delay_1239___cond_957;
  reg signed [8-1:0] __delay_data_1259__delay_1258__delay_1257__delay_1256___cond_964;
  reg [8-1:0] __delay_data_1276__delay_1275__delay_1274___plus_1025;
  reg [1-1:0] __delay_data_1294__delay_1293__delay_1292__delay_1291___eq_1031;
  reg [1-1:0] __delay_data_1323__delay_1322__delay_1321__delay_1320___eq_1034;
  reg signed [32-1:0] __delay_data_1243__delay_1242__delay_1241__delay_1240___cond_957;
  reg signed [8-1:0] __delay_data_1260__delay_1259__delay_1258__delay_1257___cond_964;
  reg [8-1:0] __delay_data_1277__delay_1276__delay_1275___plus_1025;
  reg [1-1:0] __delay_data_1295__delay_1294__delay_1293__delay_1292___eq_1031;
  reg [1-1:0] __delay_data_1324__delay_1323__delay_1322__delay_1321___eq_1034;
  wire signed [32-1:0] __substreamoutput_data_1021;
  assign __substreamoutput_data_1021 = acc_1_sum_data;
  wire [1-1:0] __substreamoutput_data_1022;
  assign __substreamoutput_data_1022 = acc_1_valid_data;
  reg signed [32-1:0] _plus_data_1023;
  reg signed [8-1:0] __delay_data_1261__delay_1260__delay_1259__delay_1258___cond_964;
  reg [8-1:0] __delay_data_1278__delay_1277__delay_1276___plus_1025;
  reg [1-1:0] __delay_data_1296__delay_1295__delay_1294__delay_1293___eq_1031;
  reg [1-1:0] __delay_data_1325__delay_1324__delay_1323__delay_1322___eq_1034;
  reg [1-1:0] __delay_data_1337__substreamoutput_1022;
  assign _mul_rshift_round_clip_4_is_root = ((_stream_matmul_55_busy)? 0 : 1) && (((_stream_conv2d_24_busy)? 0 : 1) && 1);
  assign _mul_rshift_round_clip_4_stream_oready = ((_stream_matmul_55_busy)? _stream_matmul_55_stream_oready : 1) && (((_stream_conv2d_24_busy)? _stream_conv2d_24_stream_oready : 1) && _mul_rshift_round_clip_4_stream_internal_oready);
  assign _stream_matmul_55_stream_internal_oready = ((_stream_matmul_55_busy)? _mul_rshift_round_clip_4_stream_internal_oready : 1) && (((_stream_matmul_55_busy)? _acc_1_stream_internal_oready : 1) && (((_stream_matmul_55_busy)? _add_tree_2_stream_internal_oready : 1) && (((_stream_matmul_55_busy)? _mul_5_stream_internal_oready : 1) && 1)));
  reg [1-1:0] __delay_data_1297__delay_1296__delay_1295__delay_1294___eq_1031;
  reg [1-1:0] __delay_data_1326__delay_1325__delay_1324__delay_1323___eq_1034;
  reg [1-1:0] __delay_data_1338__delay_1337__substreamoutput_1022;
  reg [1-1:0] __delay_data_1298__delay_1297__delay_1296__delay_1295___eq_1031;
  reg [1-1:0] __delay_data_1327__delay_1326__delay_1325__delay_1324___eq_1034;
  reg [1-1:0] __delay_data_1339__delay_1338____substreamoutput_1022;
  reg [1-1:0] __delay_data_1299__delay_1298__delay_1297__delay_1296___eq_1031;
  reg [1-1:0] __delay_data_1328__delay_1327__delay_1326__delay_1325___eq_1034;
  reg [1-1:0] __delay_data_1340__delay_1339____substreamoutput_1022;
  reg [1-1:0] __delay_data_1300__delay_1299__delay_1298__delay_1297___eq_1031;
  reg [1-1:0] __delay_data_1329__delay_1328__delay_1327__delay_1326___eq_1034;
  reg [1-1:0] __delay_data_1341__delay_1340____substreamoutput_1022;
  reg [1-1:0] __delay_data_1301__delay_1300__delay_1299__delay_1298___eq_1031;
  reg [1-1:0] __delay_data_1330__delay_1329__delay_1328__delay_1327___eq_1034;
  reg [1-1:0] __delay_data_1342__delay_1341____substreamoutput_1022;
  reg [1-1:0] __delay_data_1302__delay_1301__delay_1300__delay_1299___eq_1031;
  reg [1-1:0] __delay_data_1331__delay_1330__delay_1329__delay_1328___eq_1034;
  reg [1-1:0] __delay_data_1343__delay_1342____substreamoutput_1022;
  reg [1-1:0] __delay_data_1303__delay_1302__delay_1301__delay_1300___eq_1031;
  reg [1-1:0] __delay_data_1332__delay_1331__delay_1330__delay_1329___eq_1034;
  reg [1-1:0] __delay_data_1344__delay_1343____substreamoutput_1022;
  reg [1-1:0] __delay_data_1304__delay_1303__delay_1302__delay_1301___eq_1031;
  reg [1-1:0] __delay_data_1333__delay_1332__delay_1331__delay_1330___eq_1034;
  reg [1-1:0] __delay_data_1345__delay_1344____substreamoutput_1022;
  reg [1-1:0] __delay_data_1305__delay_1304__delay_1303__delay_1302___eq_1031;
  reg [1-1:0] __delay_data_1334__delay_1333__delay_1332__delay_1331___eq_1034;
  reg [1-1:0] __delay_data_1346__delay_1345____substreamoutput_1022;
  wire signed [8-1:0] __substreamoutput_data_1026;
  assign __substreamoutput_data_1026 = mul_rshift_round_clip_4_z_data;
  reg [1-1:0] _greaterthan_data_1028;
  reg signed [8-1:0] __delay_data_1279__substreamoutput_1026;
  reg [1-1:0] __delay_data_1306__delay_1305__delay_1304__delay_1303___eq_1031;
  reg [1-1:0] __delay_data_1335__delay_1334__delay_1333__delay_1332___eq_1034;
  reg [1-1:0] __delay_data_1347__delay_1346____substreamoutput_1022;
  reg signed [8-1:0] _cond_data_1030;
  reg [1-1:0] __delay_data_1307__delay_1306__delay_1305__delay_1304___eq_1031;
  reg signed [8-1:0] __delay_data_1308__delay_1279__substreamoutput_1026;
  reg [1-1:0] __delay_data_1336__delay_1335__delay_1334__delay_1333___eq_1034;
  reg [1-1:0] __delay_data_1348__delay_1347____substreamoutput_1022;
  wire signed [8-1:0] _cond_data_1033;
  assign _cond_data_1033 = (__delay_data_1307__delay_1306__delay_1305__delay_1304___eq_1031)? _cond_data_1030 : __delay_data_1308__delay_1279__substreamoutput_1026;
  wire signed [8-1:0] _cond_data_1036;
  assign _cond_data_1036 = (__delay_data_1336__delay_1335__delay_1334__delay_1333___eq_1034)? __delay_data_1308__delay_1279__substreamoutput_1026 : _cond_data_1033;
  wire signed [8-1:0] _reinterpretcast_src_1037;
  assign _reinterpretcast_src_1037 = _cond_data_1036;
  wire signed [8-1:0] _reinterpretcast_data_1037;
  assign _reinterpretcast_data_1037 = _reinterpretcast_src_1037;
  wire signed [8-1:0] stream_matmul_55_sink_26_data;
  assign stream_matmul_55_sink_26_data = _reinterpretcast_data_1037;
  wire [1-1:0] stream_matmul_55_sink_27_data;
  assign stream_matmul_55_sink_27_data = __delay_data_1348__delay_1347____substreamoutput_1022;
  wire _set_flag_1656;
  assign _set_flag_1656 = matmul_55_comp_fsm == 3;
  reg [15-1:0] __variable_wdata_936;
  assign stream_matmul_55_parameter_0_data = __variable_wdata_936;
  wire _set_flag_1657;
  assign _set_flag_1657 = matmul_55_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_937;
  assign stream_matmul_55_parameter_1_data = __variable_wdata_937;
  wire _set_flag_1658;
  assign _set_flag_1658 = matmul_55_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_938;
  assign stream_matmul_55_parameter_2_data = __variable_wdata_938;
  wire _set_flag_1659;
  assign _set_flag_1659 = matmul_55_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_939;
  assign stream_matmul_55_parameter_3_data = __variable_wdata_939;
  wire _set_flag_1660;
  assign _set_flag_1660 = matmul_55_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_940;
  assign stream_matmul_55_parameter_4_data = __variable_wdata_940;
  wire _set_flag_1661;
  assign _set_flag_1661 = matmul_55_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_951;
  assign stream_matmul_55_parameter_6_data = __variable_wdata_951;
  reg [32-1:0] _source_stream_matmul_55_source_7_pat_cur_offset_0;
  reg [32-1:0] _source_stream_matmul_55_source_7_pat_cur_offset_1;
  reg [32-1:0] _source_stream_matmul_55_source_7_pat_cur_offset_2;
  reg [32-1:0] _source_stream_matmul_55_source_7_pat_cur_offset_3;
  reg [33-1:0] _source_stream_matmul_55_source_7_pat_size_0;
  reg [33-1:0] _source_stream_matmul_55_source_7_pat_size_1;
  reg [33-1:0] _source_stream_matmul_55_source_7_pat_size_2;
  reg [33-1:0] _source_stream_matmul_55_source_7_pat_size_3;
  reg [32-1:0] _source_stream_matmul_55_source_7_pat_stride_0;
  reg [32-1:0] _source_stream_matmul_55_source_7_pat_stride_1;
  reg [32-1:0] _source_stream_matmul_55_source_7_pat_stride_2;
  reg [32-1:0] _source_stream_matmul_55_source_7_pat_stride_3;
  reg [33-1:0] _source_stream_matmul_55_source_7_pat_count_0;
  reg [33-1:0] _source_stream_matmul_55_source_7_pat_count_1;
  reg [33-1:0] _source_stream_matmul_55_source_7_pat_count_2;
  reg [33-1:0] _source_stream_matmul_55_source_7_pat_count_3;
  reg [33-1:0] _source_stream_matmul_55_source_7_pat_size_buf_0;
  reg [33-1:0] _source_stream_matmul_55_source_7_pat_size_buf_1;
  reg [33-1:0] _source_stream_matmul_55_source_7_pat_size_buf_2;
  reg [33-1:0] _source_stream_matmul_55_source_7_pat_size_buf_3;
  reg [32-1:0] _source_stream_matmul_55_source_7_pat_stride_buf_0;
  reg [32-1:0] _source_stream_matmul_55_source_7_pat_stride_buf_1;
  reg [32-1:0] _source_stream_matmul_55_source_7_pat_stride_buf_2;
  reg [32-1:0] _source_stream_matmul_55_source_7_pat_stride_buf_3;
  wire _set_flag_1662;
  assign _set_flag_1662 = matmul_55_comp_fsm == 3;
  assign ram_w32_l4096_id0_0_addr = (_stream_matmul_55_stream_oready && _stream_matmul_55_source_7_source_ram_renable && (_stream_matmul_55_source_7_source_sel == 1))? _stream_matmul_55_source_7_source_ram_raddr : 
                                    (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_7_source_ram_renable && (_stream_conv2d_24_source_7_source_sel == 1))? _stream_conv2d_24_source_7_source_ram_raddr : 'hx;
  assign ram_w32_l4096_id0_0_enable = (_stream_matmul_55_stream_oready && _stream_matmul_55_source_7_source_ram_renable && (_stream_matmul_55_source_7_source_sel == 1))? 1'd1 : 
                                      (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_7_source_ram_renable && (_stream_conv2d_24_source_7_source_sel == 1))? 1'd1 : 0;
  localparam _tmp_1663 = 1;
  wire [_tmp_1663-1:0] _tmp_1664;
  assign _tmp_1664 = _stream_matmul_55_stream_oready && _stream_matmul_55_source_7_source_ram_renable && (_stream_matmul_55_source_7_source_sel == 1);
  reg [_tmp_1663-1:0] __tmp_1664_1;
  assign _stream_matmul_55_source_7_source_ram_rdata = (_stream_matmul_55_source_7_source_sel == 1)? ram_w32_l4096_id0_0_rdata : 'hx;
  reg [32-1:0] __variable_wdata_952;
  assign stream_matmul_55_source_7_data = __variable_wdata_952;
  reg [32-1:0] _stream_matmul_55_source_7_source_pat_fsm_0;
  localparam _stream_matmul_55_source_7_source_pat_fsm_0_init = 0;
  wire [32-1:0] _stream_matmul_55_source_7_source_pat_all_offset;
  assign _stream_matmul_55_source_7_source_pat_all_offset = _stream_matmul_55_source_7_source_offset_buf + _source_stream_matmul_55_source_7_pat_cur_offset_0 + _source_stream_matmul_55_source_7_pat_cur_offset_1 + _source_stream_matmul_55_source_7_pat_cur_offset_2 + _source_stream_matmul_55_source_7_pat_cur_offset_3;
  wire _set_flag_1665;
  assign _set_flag_1665 = matmul_55_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_958;
  assign stream_matmul_55_parameter_8_data = __variable_wdata_958;
  reg [32-1:0] _source_stream_matmul_55_source_9_pat_cur_offset_0;
  reg [32-1:0] _source_stream_matmul_55_source_9_pat_cur_offset_1;
  reg [32-1:0] _source_stream_matmul_55_source_9_pat_cur_offset_2;
  reg [32-1:0] _source_stream_matmul_55_source_9_pat_cur_offset_3;
  reg [33-1:0] _source_stream_matmul_55_source_9_pat_size_0;
  reg [33-1:0] _source_stream_matmul_55_source_9_pat_size_1;
  reg [33-1:0] _source_stream_matmul_55_source_9_pat_size_2;
  reg [33-1:0] _source_stream_matmul_55_source_9_pat_size_3;
  reg [32-1:0] _source_stream_matmul_55_source_9_pat_stride_0;
  reg [32-1:0] _source_stream_matmul_55_source_9_pat_stride_1;
  reg [32-1:0] _source_stream_matmul_55_source_9_pat_stride_2;
  reg [32-1:0] _source_stream_matmul_55_source_9_pat_stride_3;
  reg [33-1:0] _source_stream_matmul_55_source_9_pat_count_0;
  reg [33-1:0] _source_stream_matmul_55_source_9_pat_count_1;
  reg [33-1:0] _source_stream_matmul_55_source_9_pat_count_2;
  reg [33-1:0] _source_stream_matmul_55_source_9_pat_count_3;
  reg [33-1:0] _source_stream_matmul_55_source_9_pat_size_buf_0;
  reg [33-1:0] _source_stream_matmul_55_source_9_pat_size_buf_1;
  reg [33-1:0] _source_stream_matmul_55_source_9_pat_size_buf_2;
  reg [33-1:0] _source_stream_matmul_55_source_9_pat_size_buf_3;
  reg [32-1:0] _source_stream_matmul_55_source_9_pat_stride_buf_0;
  reg [32-1:0] _source_stream_matmul_55_source_9_pat_stride_buf_1;
  reg [32-1:0] _source_stream_matmul_55_source_9_pat_stride_buf_2;
  reg [32-1:0] _source_stream_matmul_55_source_9_pat_stride_buf_3;
  wire _set_flag_1666;
  assign _set_flag_1666 = matmul_55_comp_fsm == 3;
  wire [2-1:0] read_rtl_bank_1667;
  assign read_rtl_bank_1667 = _stream_matmul_55_source_9_source_ram_raddr;
  reg [2-1:0] _tmp_1668;
  assign ram_w8_l2048_id0_0_0_addr = (_stream_matmul_55_stream_oready && _stream_matmul_55_source_9_source_ram_renable && (_stream_matmul_55_source_9_source_sel == 2))? _stream_matmul_55_source_9_source_ram_raddr >> 2 : 
                                     (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_9_source_ram_renable && (_stream_conv2d_24_source_9_source_sel == 2))? _stream_conv2d_24_source_9_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l2048_id0_0_0_enable = (_stream_matmul_55_stream_oready && _stream_matmul_55_source_9_source_ram_renable && (_stream_matmul_55_source_9_source_sel == 2))? 1'd1 : 
                                       (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_9_source_ram_renable && (_stream_conv2d_24_source_9_source_sel == 2))? 1'd1 : 0;
  localparam _tmp_1669 = 1;
  wire [_tmp_1669-1:0] _tmp_1670;
  assign _tmp_1670 = _stream_matmul_55_stream_oready && _stream_matmul_55_source_9_source_ram_renable && (_stream_matmul_55_source_9_source_sel == 2);
  reg [_tmp_1669-1:0] __tmp_1670_1;
  assign ram_w8_l2048_id0_1_0_addr = (_stream_matmul_55_stream_oready && _stream_matmul_55_source_9_source_ram_renable && (_stream_matmul_55_source_9_source_sel == 2))? _stream_matmul_55_source_9_source_ram_raddr >> 2 : 
                                     (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_9_source_ram_renable && (_stream_conv2d_24_source_9_source_sel == 2))? _stream_conv2d_24_source_9_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l2048_id0_1_0_enable = (_stream_matmul_55_stream_oready && _stream_matmul_55_source_9_source_ram_renable && (_stream_matmul_55_source_9_source_sel == 2))? 1'd1 : 
                                       (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_9_source_ram_renable && (_stream_conv2d_24_source_9_source_sel == 2))? 1'd1 : 0;
  localparam _tmp_1671 = 1;
  wire [_tmp_1671-1:0] _tmp_1672;
  assign _tmp_1672 = _stream_matmul_55_stream_oready && _stream_matmul_55_source_9_source_ram_renable && (_stream_matmul_55_source_9_source_sel == 2);
  reg [_tmp_1671-1:0] __tmp_1672_1;
  assign ram_w8_l2048_id0_2_0_addr = (_stream_matmul_55_stream_oready && _stream_matmul_55_source_9_source_ram_renable && (_stream_matmul_55_source_9_source_sel == 2))? _stream_matmul_55_source_9_source_ram_raddr >> 2 : 
                                     (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_9_source_ram_renable && (_stream_conv2d_24_source_9_source_sel == 2))? _stream_conv2d_24_source_9_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l2048_id0_2_0_enable = (_stream_matmul_55_stream_oready && _stream_matmul_55_source_9_source_ram_renable && (_stream_matmul_55_source_9_source_sel == 2))? 1'd1 : 
                                       (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_9_source_ram_renable && (_stream_conv2d_24_source_9_source_sel == 2))? 1'd1 : 0;
  localparam _tmp_1673 = 1;
  wire [_tmp_1673-1:0] _tmp_1674;
  assign _tmp_1674 = _stream_matmul_55_stream_oready && _stream_matmul_55_source_9_source_ram_renable && (_stream_matmul_55_source_9_source_sel == 2);
  reg [_tmp_1673-1:0] __tmp_1674_1;
  assign ram_w8_l2048_id0_3_0_addr = (_stream_matmul_55_stream_oready && _stream_matmul_55_source_9_source_ram_renable && (_stream_matmul_55_source_9_source_sel == 2))? _stream_matmul_55_source_9_source_ram_raddr >> 2 : 
                                     (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_9_source_ram_renable && (_stream_conv2d_24_source_9_source_sel == 2))? _stream_conv2d_24_source_9_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l2048_id0_3_0_enable = (_stream_matmul_55_stream_oready && _stream_matmul_55_source_9_source_ram_renable && (_stream_matmul_55_source_9_source_sel == 2))? 1'd1 : 
                                       (_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_9_source_ram_renable && (_stream_conv2d_24_source_9_source_sel == 2))? 1'd1 : 0;
  localparam _tmp_1675 = 1;
  wire [_tmp_1675-1:0] _tmp_1676;
  assign _tmp_1676 = _stream_matmul_55_stream_oready && _stream_matmul_55_source_9_source_ram_renable && (_stream_matmul_55_source_9_source_sel == 2);
  reg [_tmp_1675-1:0] __tmp_1676_1;
  wire signed [8-1:0] read_rtl_rdata_1677;
  wire read_rtl_rvalid_1678;
  assign read_rtl_rdata_1677 = (_tmp_1668 == 0)? ram_w8_l2048_id0_0_0_rdata : 
                               (_tmp_1668 == 1)? ram_w8_l2048_id0_1_0_rdata : 
                               (_tmp_1668 == 2)? ram_w8_l2048_id0_2_0_rdata : 
                               (_tmp_1668 == 3)? ram_w8_l2048_id0_3_0_rdata : 0;
  assign read_rtl_rvalid_1678 = __tmp_1670_1;
  assign _stream_matmul_55_source_9_source_ram_rdata = (_stream_matmul_55_source_9_source_sel == 2)? read_rtl_rdata_1677 : 'hx;
  reg [8-1:0] __variable_wdata_959;
  assign stream_matmul_55_source_9_data = __variable_wdata_959;
  reg [32-1:0] _stream_matmul_55_source_9_source_pat_fsm_1;
  localparam _stream_matmul_55_source_9_source_pat_fsm_1_init = 0;
  wire [32-1:0] _stream_matmul_55_source_9_source_pat_all_offset;
  assign _stream_matmul_55_source_9_source_pat_all_offset = _stream_matmul_55_source_9_source_offset_buf + _source_stream_matmul_55_source_9_pat_cur_offset_0 + _source_stream_matmul_55_source_9_pat_cur_offset_1 + _source_stream_matmul_55_source_9_pat_cur_offset_2 + _source_stream_matmul_55_source_9_pat_cur_offset_3;
  wire _set_flag_1679;
  assign _set_flag_1679 = matmul_55_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_965;
  assign stream_matmul_55_parameter_10_data = __variable_wdata_965;
  wire _set_flag_1680;
  assign _set_flag_1680 = matmul_55_comp_fsm == 3;
  reg [8-1:0] __variable_wdata_966;
  assign stream_matmul_55_source_11_data = __variable_wdata_966;
  wire _set_flag_1681;
  assign _set_flag_1681 = matmul_55_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_972;
  assign stream_matmul_55_parameter_12_data = __variable_wdata_972;
  wire _set_flag_1682;
  assign _set_flag_1682 = matmul_55_comp_fsm == 3;
  reg [8-1:0] __variable_wdata_973;
  assign stream_matmul_55_source_13_data = __variable_wdata_973;
  wire _set_flag_1683;
  assign _set_flag_1683 = matmul_55_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_979;
  assign stream_matmul_55_parameter_14_data = __variable_wdata_979;
  wire _set_flag_1684;
  assign _set_flag_1684 = matmul_55_comp_fsm == 3;
  reg [8-1:0] __variable_wdata_980;
  assign stream_matmul_55_source_15_data = __variable_wdata_980;
  wire _set_flag_1685;
  assign _set_flag_1685 = matmul_55_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_986;
  assign stream_matmul_55_parameter_16_data = __variable_wdata_986;
  wire _set_flag_1686;
  assign _set_flag_1686 = matmul_55_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_987;
  assign stream_matmul_55_parameter_17_data = __variable_wdata_987;
  wire _set_flag_1687;
  assign _set_flag_1687 = matmul_55_comp_fsm == 3;
  reg [5-1:0] __variable_wdata_988;
  assign stream_matmul_55_parameter_18_data = __variable_wdata_988;
  wire _set_flag_1688;
  assign _set_flag_1688 = matmul_55_comp_fsm == 3;
  reg [2-1:0] __variable_wdata_989;
  assign stream_matmul_55_parameter_19_data = __variable_wdata_989;
  reg [32-1:0] _source_stream_matmul_55_source_20_pat_cur_offset_0;
  reg [32-1:0] _source_stream_matmul_55_source_20_pat_cur_offset_1;
  reg [32-1:0] _source_stream_matmul_55_source_20_pat_cur_offset_2;
  reg [32-1:0] _source_stream_matmul_55_source_20_pat_cur_offset_3;
  reg [33-1:0] _source_stream_matmul_55_source_20_pat_size_0;
  reg [33-1:0] _source_stream_matmul_55_source_20_pat_size_1;
  reg [33-1:0] _source_stream_matmul_55_source_20_pat_size_2;
  reg [33-1:0] _source_stream_matmul_55_source_20_pat_size_3;
  reg [32-1:0] _source_stream_matmul_55_source_20_pat_stride_0;
  reg [32-1:0] _source_stream_matmul_55_source_20_pat_stride_1;
  reg [32-1:0] _source_stream_matmul_55_source_20_pat_stride_2;
  reg [32-1:0] _source_stream_matmul_55_source_20_pat_stride_3;
  reg [33-1:0] _source_stream_matmul_55_source_20_pat_count_0;
  reg [33-1:0] _source_stream_matmul_55_source_20_pat_count_1;
  reg [33-1:0] _source_stream_matmul_55_source_20_pat_count_2;
  reg [33-1:0] _source_stream_matmul_55_source_20_pat_count_3;
  reg [33-1:0] _source_stream_matmul_55_source_20_pat_size_buf_0;
  reg [33-1:0] _source_stream_matmul_55_source_20_pat_size_buf_1;
  reg [33-1:0] _source_stream_matmul_55_source_20_pat_size_buf_2;
  reg [33-1:0] _source_stream_matmul_55_source_20_pat_size_buf_3;
  reg [32-1:0] _source_stream_matmul_55_source_20_pat_stride_buf_0;
  reg [32-1:0] _source_stream_matmul_55_source_20_pat_stride_buf_1;
  reg [32-1:0] _source_stream_matmul_55_source_20_pat_stride_buf_2;
  reg [32-1:0] _source_stream_matmul_55_source_20_pat_stride_buf_3;
  wire _set_flag_1689;
  assign _set_flag_1689 = matmul_55_comp_fsm == 3;
  wire [2-1:0] read_rtl_bank_1690;
  assign read_rtl_bank_1690 = _stream_matmul_55_source_20_source_ram_raddr;
  reg [2-1:0] _tmp_1691;
  assign ram_w8_l32768_id0_0_0_addr = (_stream_matmul_55_stream_oready && _stream_matmul_55_source_20_source_ram_renable && (_stream_matmul_55_source_20_source_sel == 3))? _stream_matmul_55_source_20_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l32768_id0_0_0_enable = (_stream_matmul_55_stream_oready && _stream_matmul_55_source_20_source_ram_renable && (_stream_matmul_55_source_20_source_sel == 3))? 1'd1 : 0;
  localparam _tmp_1692 = 1;
  wire [_tmp_1692-1:0] _tmp_1693;
  assign _tmp_1693 = _stream_matmul_55_stream_oready && _stream_matmul_55_source_20_source_ram_renable && (_stream_matmul_55_source_20_source_sel == 3);
  reg [_tmp_1692-1:0] __tmp_1693_1;
  assign ram_w8_l32768_id0_1_0_addr = (_stream_matmul_55_stream_oready && _stream_matmul_55_source_20_source_ram_renable && (_stream_matmul_55_source_20_source_sel == 3))? _stream_matmul_55_source_20_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l32768_id0_1_0_enable = (_stream_matmul_55_stream_oready && _stream_matmul_55_source_20_source_ram_renable && (_stream_matmul_55_source_20_source_sel == 3))? 1'd1 : 0;
  localparam _tmp_1694 = 1;
  wire [_tmp_1694-1:0] _tmp_1695;
  assign _tmp_1695 = _stream_matmul_55_stream_oready && _stream_matmul_55_source_20_source_ram_renable && (_stream_matmul_55_source_20_source_sel == 3);
  reg [_tmp_1694-1:0] __tmp_1695_1;
  assign ram_w8_l32768_id0_2_0_addr = (_stream_matmul_55_stream_oready && _stream_matmul_55_source_20_source_ram_renable && (_stream_matmul_55_source_20_source_sel == 3))? _stream_matmul_55_source_20_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l32768_id0_2_0_enable = (_stream_matmul_55_stream_oready && _stream_matmul_55_source_20_source_ram_renable && (_stream_matmul_55_source_20_source_sel == 3))? 1'd1 : 0;
  localparam _tmp_1696 = 1;
  wire [_tmp_1696-1:0] _tmp_1697;
  assign _tmp_1697 = _stream_matmul_55_stream_oready && _stream_matmul_55_source_20_source_ram_renable && (_stream_matmul_55_source_20_source_sel == 3);
  reg [_tmp_1696-1:0] __tmp_1697_1;
  assign ram_w8_l32768_id0_3_0_addr = (_stream_matmul_55_stream_oready && _stream_matmul_55_source_20_source_ram_renable && (_stream_matmul_55_source_20_source_sel == 3))? _stream_matmul_55_source_20_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l32768_id0_3_0_enable = (_stream_matmul_55_stream_oready && _stream_matmul_55_source_20_source_ram_renable && (_stream_matmul_55_source_20_source_sel == 3))? 1'd1 : 0;
  localparam _tmp_1698 = 1;
  wire [_tmp_1698-1:0] _tmp_1699;
  assign _tmp_1699 = _stream_matmul_55_stream_oready && _stream_matmul_55_source_20_source_ram_renable && (_stream_matmul_55_source_20_source_sel == 3);
  reg [_tmp_1698-1:0] __tmp_1699_1;
  wire signed [8-1:0] read_rtl_rdata_1700;
  wire read_rtl_rvalid_1701;
  assign read_rtl_rdata_1700 = (_tmp_1691 == 0)? ram_w8_l32768_id0_0_0_rdata : 
                               (_tmp_1691 == 1)? ram_w8_l32768_id0_1_0_rdata : 
                               (_tmp_1691 == 2)? ram_w8_l32768_id0_2_0_rdata : 
                               (_tmp_1691 == 3)? ram_w8_l32768_id0_3_0_rdata : 0;
  assign read_rtl_rvalid_1701 = __tmp_1693_1;
  assign _stream_matmul_55_source_20_source_ram_rdata = (_stream_matmul_55_source_20_source_sel == 3)? read_rtl_rdata_1700 : 'hx;
  reg [8-1:0] __variable_wdata_990;
  assign stream_matmul_55_source_20_data = __variable_wdata_990;
  reg [32-1:0] _stream_matmul_55_source_20_source_pat_fsm_2;
  localparam _stream_matmul_55_source_20_source_pat_fsm_2_init = 0;
  wire [32-1:0] _stream_matmul_55_source_20_source_pat_all_offset;
  assign _stream_matmul_55_source_20_source_pat_all_offset = _stream_matmul_55_source_20_source_offset_buf + _source_stream_matmul_55_source_20_pat_cur_offset_0 + _source_stream_matmul_55_source_20_pat_cur_offset_1 + _source_stream_matmul_55_source_20_pat_cur_offset_2 + _source_stream_matmul_55_source_20_pat_cur_offset_3;
  reg [32-1:0] _source_stream_matmul_55_source_21_pat_cur_offset_0;
  reg [32-1:0] _source_stream_matmul_55_source_21_pat_cur_offset_1;
  reg [32-1:0] _source_stream_matmul_55_source_21_pat_cur_offset_2;
  reg [32-1:0] _source_stream_matmul_55_source_21_pat_cur_offset_3;
  reg [33-1:0] _source_stream_matmul_55_source_21_pat_size_0;
  reg [33-1:0] _source_stream_matmul_55_source_21_pat_size_1;
  reg [33-1:0] _source_stream_matmul_55_source_21_pat_size_2;
  reg [33-1:0] _source_stream_matmul_55_source_21_pat_size_3;
  reg [32-1:0] _source_stream_matmul_55_source_21_pat_stride_0;
  reg [32-1:0] _source_stream_matmul_55_source_21_pat_stride_1;
  reg [32-1:0] _source_stream_matmul_55_source_21_pat_stride_2;
  reg [32-1:0] _source_stream_matmul_55_source_21_pat_stride_3;
  reg [33-1:0] _source_stream_matmul_55_source_21_pat_count_0;
  reg [33-1:0] _source_stream_matmul_55_source_21_pat_count_1;
  reg [33-1:0] _source_stream_matmul_55_source_21_pat_count_2;
  reg [33-1:0] _source_stream_matmul_55_source_21_pat_count_3;
  reg [33-1:0] _source_stream_matmul_55_source_21_pat_size_buf_0;
  reg [33-1:0] _source_stream_matmul_55_source_21_pat_size_buf_1;
  reg [33-1:0] _source_stream_matmul_55_source_21_pat_size_buf_2;
  reg [33-1:0] _source_stream_matmul_55_source_21_pat_size_buf_3;
  reg [32-1:0] _source_stream_matmul_55_source_21_pat_stride_buf_0;
  reg [32-1:0] _source_stream_matmul_55_source_21_pat_stride_buf_1;
  reg [32-1:0] _source_stream_matmul_55_source_21_pat_stride_buf_2;
  reg [32-1:0] _source_stream_matmul_55_source_21_pat_stride_buf_3;
  wire _set_flag_1702;
  assign _set_flag_1702 = matmul_55_comp_fsm == 3;
  wire [2-1:0] read_rtl_bank_1703;
  assign read_rtl_bank_1703 = _stream_matmul_55_source_21_source_ram_raddr;
  reg [2-1:0] _tmp_1704;
  assign ram_w8_l262144_id0_0_0_addr = (_stream_matmul_55_stream_oready && _stream_matmul_55_source_21_source_ram_renable && (_stream_matmul_55_source_21_source_sel == 4))? _stream_matmul_55_source_21_source_ram_raddr >> 2 : 
                                       (_stream_max_pool_serial_26_stream_oready && _stream_max_pool_serial_26_source_1_source_ram_renable && (_stream_max_pool_serial_26_source_1_source_sel == 1))? _stream_max_pool_serial_26_source_1_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l262144_id0_0_0_enable = (_stream_matmul_55_stream_oready && _stream_matmul_55_source_21_source_ram_renable && (_stream_matmul_55_source_21_source_sel == 4))? 1'd1 : 
                                         (_stream_max_pool_serial_26_stream_oready && _stream_max_pool_serial_26_source_1_source_ram_renable && (_stream_max_pool_serial_26_source_1_source_sel == 1))? 1'd1 : 0;
  localparam _tmp_1705 = 1;
  wire [_tmp_1705-1:0] _tmp_1706;
  assign _tmp_1706 = _stream_matmul_55_stream_oready && _stream_matmul_55_source_21_source_ram_renable && (_stream_matmul_55_source_21_source_sel == 4);
  reg [_tmp_1705-1:0] __tmp_1706_1;
  assign ram_w8_l262144_id0_1_0_addr = (_stream_matmul_55_stream_oready && _stream_matmul_55_source_21_source_ram_renable && (_stream_matmul_55_source_21_source_sel == 4))? _stream_matmul_55_source_21_source_ram_raddr >> 2 : 
                                       (_stream_max_pool_serial_26_stream_oready && _stream_max_pool_serial_26_source_1_source_ram_renable && (_stream_max_pool_serial_26_source_1_source_sel == 1))? _stream_max_pool_serial_26_source_1_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l262144_id0_1_0_enable = (_stream_matmul_55_stream_oready && _stream_matmul_55_source_21_source_ram_renable && (_stream_matmul_55_source_21_source_sel == 4))? 1'd1 : 
                                         (_stream_max_pool_serial_26_stream_oready && _stream_max_pool_serial_26_source_1_source_ram_renable && (_stream_max_pool_serial_26_source_1_source_sel == 1))? 1'd1 : 0;
  localparam _tmp_1707 = 1;
  wire [_tmp_1707-1:0] _tmp_1708;
  assign _tmp_1708 = _stream_matmul_55_stream_oready && _stream_matmul_55_source_21_source_ram_renable && (_stream_matmul_55_source_21_source_sel == 4);
  reg [_tmp_1707-1:0] __tmp_1708_1;
  assign ram_w8_l262144_id0_2_0_addr = (_stream_matmul_55_stream_oready && _stream_matmul_55_source_21_source_ram_renable && (_stream_matmul_55_source_21_source_sel == 4))? _stream_matmul_55_source_21_source_ram_raddr >> 2 : 
                                       (_stream_max_pool_serial_26_stream_oready && _stream_max_pool_serial_26_source_1_source_ram_renable && (_stream_max_pool_serial_26_source_1_source_sel == 1))? _stream_max_pool_serial_26_source_1_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l262144_id0_2_0_enable = (_stream_matmul_55_stream_oready && _stream_matmul_55_source_21_source_ram_renable && (_stream_matmul_55_source_21_source_sel == 4))? 1'd1 : 
                                         (_stream_max_pool_serial_26_stream_oready && _stream_max_pool_serial_26_source_1_source_ram_renable && (_stream_max_pool_serial_26_source_1_source_sel == 1))? 1'd1 : 0;
  localparam _tmp_1709 = 1;
  wire [_tmp_1709-1:0] _tmp_1710;
  assign _tmp_1710 = _stream_matmul_55_stream_oready && _stream_matmul_55_source_21_source_ram_renable && (_stream_matmul_55_source_21_source_sel == 4);
  reg [_tmp_1709-1:0] __tmp_1710_1;
  assign ram_w8_l262144_id0_3_0_addr = (_stream_matmul_55_stream_oready && _stream_matmul_55_source_21_source_ram_renable && (_stream_matmul_55_source_21_source_sel == 4))? _stream_matmul_55_source_21_source_ram_raddr >> 2 : 
                                       (_stream_max_pool_serial_26_stream_oready && _stream_max_pool_serial_26_source_1_source_ram_renable && (_stream_max_pool_serial_26_source_1_source_sel == 1))? _stream_max_pool_serial_26_source_1_source_ram_raddr >> 2 : 'hx;
  assign ram_w8_l262144_id0_3_0_enable = (_stream_matmul_55_stream_oready && _stream_matmul_55_source_21_source_ram_renable && (_stream_matmul_55_source_21_source_sel == 4))? 1'd1 : 
                                         (_stream_max_pool_serial_26_stream_oready && _stream_max_pool_serial_26_source_1_source_ram_renable && (_stream_max_pool_serial_26_source_1_source_sel == 1))? 1'd1 : 0;
  localparam _tmp_1711 = 1;
  wire [_tmp_1711-1:0] _tmp_1712;
  assign _tmp_1712 = _stream_matmul_55_stream_oready && _stream_matmul_55_source_21_source_ram_renable && (_stream_matmul_55_source_21_source_sel == 4);
  reg [_tmp_1711-1:0] __tmp_1712_1;
  wire signed [8-1:0] read_rtl_rdata_1713;
  wire read_rtl_rvalid_1714;
  assign read_rtl_rdata_1713 = (_tmp_1704 == 0)? ram_w8_l262144_id0_0_0_rdata : 
                               (_tmp_1704 == 1)? ram_w8_l262144_id0_1_0_rdata : 
                               (_tmp_1704 == 2)? ram_w8_l262144_id0_2_0_rdata : 
                               (_tmp_1704 == 3)? ram_w8_l262144_id0_3_0_rdata : 0;
  assign read_rtl_rvalid_1714 = __tmp_1706_1;
  assign _stream_matmul_55_source_21_source_ram_rdata = (_stream_matmul_55_source_21_source_sel == 4)? read_rtl_rdata_1713 : 'hx;
  reg [8-1:0] __variable_wdata_1004;
  assign stream_matmul_55_source_21_data = __variable_wdata_1004;
  reg [32-1:0] _stream_matmul_55_source_21_source_pat_fsm_3;
  localparam _stream_matmul_55_source_21_source_pat_fsm_3_init = 0;
  wire [32-1:0] _stream_matmul_55_source_21_source_pat_all_offset;
  assign _stream_matmul_55_source_21_source_pat_all_offset = _stream_matmul_55_source_21_source_offset_buf + _source_stream_matmul_55_source_21_pat_cur_offset_0 + _source_stream_matmul_55_source_21_pat_cur_offset_1 + _source_stream_matmul_55_source_21_pat_cur_offset_2 + _source_stream_matmul_55_source_21_pat_cur_offset_3;
  wire _set_flag_1715;
  assign _set_flag_1715 = matmul_55_comp_fsm == 3;
  reg _tmp_1716;
  reg _tmp_1717;
  reg _tmp_1718;
  reg _tmp_1719;
  reg _tmp_1720;
  reg _tmp_1721;
  reg _tmp_1722;
  reg _tmp_1723;
  reg _tmp_1724;
  reg _tmp_1725;
  reg _tmp_1726;
  reg _tmp_1727;
  reg _tmp_1728;
  reg _tmp_1729;
  reg _tmp_1730;
  reg _tmp_1731;
  reg _tmp_1732;
  reg _tmp_1733;
  reg _tmp_1734;
  reg _tmp_1735;
  reg _tmp_1736;
  reg _tmp_1737;
  reg _tmp_1738;
  reg _tmp_1739;
  reg _tmp_1740;
  reg _tmp_1741;
  reg _tmp_1742;
  reg _tmp_1743;
  reg _tmp_1744;
  reg _tmp_1745;
  reg _tmp_1746;
  localparam _tmp_1747 = 33;
  wire [_tmp_1747-1:0] _tmp_1748;
  assign _tmp_1748 = matmul_55_stream_out_local + matmul_55_out_page_comp_offset_buf;
  reg [_tmp_1747-1:0] _tmp_1749;
  reg [_tmp_1747-1:0] _tmp_1750;
  reg [_tmp_1747-1:0] _tmp_1751;
  reg [_tmp_1747-1:0] _tmp_1752;
  reg [_tmp_1747-1:0] _tmp_1753;
  reg [_tmp_1747-1:0] _tmp_1754;
  reg [_tmp_1747-1:0] _tmp_1755;
  reg [_tmp_1747-1:0] _tmp_1756;
  reg [_tmp_1747-1:0] _tmp_1757;
  reg [_tmp_1747-1:0] _tmp_1758;
  reg [_tmp_1747-1:0] _tmp_1759;
  reg [_tmp_1747-1:0] _tmp_1760;
  reg [_tmp_1747-1:0] _tmp_1761;
  reg [_tmp_1747-1:0] _tmp_1762;
  reg [_tmp_1747-1:0] _tmp_1763;
  reg [_tmp_1747-1:0] _tmp_1764;
  reg [_tmp_1747-1:0] _tmp_1765;
  reg [_tmp_1747-1:0] _tmp_1766;
  reg [_tmp_1747-1:0] _tmp_1767;
  reg [_tmp_1747-1:0] _tmp_1768;
  reg [_tmp_1747-1:0] _tmp_1769;
  reg [_tmp_1747-1:0] _tmp_1770;
  reg [_tmp_1747-1:0] _tmp_1771;
  reg [_tmp_1747-1:0] _tmp_1772;
  reg [_tmp_1747-1:0] _tmp_1773;
  reg [_tmp_1747-1:0] _tmp_1774;
  reg [_tmp_1747-1:0] _tmp_1775;
  reg [_tmp_1747-1:0] _tmp_1776;
  reg [_tmp_1747-1:0] _tmp_1777;
  reg [_tmp_1747-1:0] _tmp_1778;
  reg [_tmp_1747-1:0] _tmp_1779;
  reg [32-1:0] _tmp_1780;
  reg [32-1:0] _tmp_1781;
  reg [32-1:0] _tmp_1782;
  reg [32-1:0] _tmp_1783;
  reg [32-1:0] _tmp_1784;
  reg [32-1:0] _tmp_1785;
  reg [32-1:0] _tmp_1786;
  reg [32-1:0] _tmp_1787;
  reg [32-1:0] _tmp_1788;
  reg [32-1:0] _tmp_1789;
  reg [32-1:0] _tmp_1790;
  reg [32-1:0] _tmp_1791;
  reg [32-1:0] _tmp_1792;
  reg [32-1:0] _tmp_1793;
  reg [32-1:0] _tmp_1794;
  reg [32-1:0] _tmp_1795;
  reg [32-1:0] _tmp_1796;
  reg [32-1:0] _tmp_1797;
  reg [32-1:0] _tmp_1798;
  reg [32-1:0] _tmp_1799;
  reg [32-1:0] _tmp_1800;
  reg [32-1:0] _tmp_1801;
  reg [32-1:0] _tmp_1802;
  reg [32-1:0] _tmp_1803;
  reg [32-1:0] _tmp_1804;
  reg [32-1:0] _tmp_1805;
  reg [32-1:0] _tmp_1806;
  reg [32-1:0] _tmp_1807;
  reg [32-1:0] _tmp_1808;
  reg [32-1:0] _tmp_1809;
  reg [32-1:0] _tmp_1810;
  wire [2-1:0] write_rtl_bank_1811;
  assign write_rtl_bank_1811 = _stream_matmul_55_sink_26_sink_waddr;
  assign ram_w8_l2048_id1_0_0_addr = (_stream_matmul_55_stream_oready && _stream_matmul_55_sink_26_sink_wenable && (_stream_matmul_55_sink_26_sink_sel == 5) && (write_rtl_bank_1811 == 0))? _stream_matmul_55_sink_26_sink_waddr >> 2 : 
                                     (_stream_conv2d_24_stream_oready && _stream_conv2d_24_sink_50_sink_wenable && (_stream_conv2d_24_sink_50_sink_sel == 21) && (write_rtl_bank_766 == 0))? _stream_conv2d_24_sink_50_sink_waddr >> 2 : 'hx;
  assign ram_w8_l2048_id1_0_0_wdata = (_stream_matmul_55_stream_oready && _stream_matmul_55_sink_26_sink_wenable && (_stream_matmul_55_sink_26_sink_sel == 5) && (write_rtl_bank_1811 == 0))? _stream_matmul_55_sink_26_sink_wdata : 
                                      (_stream_conv2d_24_stream_oready && _stream_conv2d_24_sink_50_sink_wenable && (_stream_conv2d_24_sink_50_sink_sel == 21) && (write_rtl_bank_766 == 0))? _stream_conv2d_24_sink_50_sink_wdata : 'hx;
  assign ram_w8_l2048_id1_0_0_wenable = (_stream_matmul_55_stream_oready && _stream_matmul_55_sink_26_sink_wenable && (_stream_matmul_55_sink_26_sink_sel == 5) && (write_rtl_bank_1811 == 0))? 1'd1 : 
                                        (_stream_conv2d_24_stream_oready && _stream_conv2d_24_sink_50_sink_wenable && (_stream_conv2d_24_sink_50_sink_sel == 21) && (write_rtl_bank_766 == 0))? 1'd1 : 0;
  assign ram_w8_l2048_id1_0_0_enable = (_stream_matmul_55_stream_oready && _stream_matmul_55_sink_26_sink_wenable && (_stream_matmul_55_sink_26_sink_sel == 5) && (write_rtl_bank_1811 == 0))? 1'd1 : 
                                       (_stream_conv2d_24_stream_oready && _stream_conv2d_24_sink_50_sink_wenable && (_stream_conv2d_24_sink_50_sink_sel == 21) && (write_rtl_bank_766 == 0))? 1'd1 : 0;
  assign ram_w8_l2048_id1_1_0_addr = (_stream_matmul_55_stream_oready && _stream_matmul_55_sink_26_sink_wenable && (_stream_matmul_55_sink_26_sink_sel == 5) && (write_rtl_bank_1811 == 1))? _stream_matmul_55_sink_26_sink_waddr >> 2 : 
                                     (_stream_conv2d_24_stream_oready && _stream_conv2d_24_sink_50_sink_wenable && (_stream_conv2d_24_sink_50_sink_sel == 21) && (write_rtl_bank_766 == 1))? _stream_conv2d_24_sink_50_sink_waddr >> 2 : 'hx;
  assign ram_w8_l2048_id1_1_0_wdata = (_stream_matmul_55_stream_oready && _stream_matmul_55_sink_26_sink_wenable && (_stream_matmul_55_sink_26_sink_sel == 5) && (write_rtl_bank_1811 == 1))? _stream_matmul_55_sink_26_sink_wdata : 
                                      (_stream_conv2d_24_stream_oready && _stream_conv2d_24_sink_50_sink_wenable && (_stream_conv2d_24_sink_50_sink_sel == 21) && (write_rtl_bank_766 == 1))? _stream_conv2d_24_sink_50_sink_wdata : 'hx;
  assign ram_w8_l2048_id1_1_0_wenable = (_stream_matmul_55_stream_oready && _stream_matmul_55_sink_26_sink_wenable && (_stream_matmul_55_sink_26_sink_sel == 5) && (write_rtl_bank_1811 == 1))? 1'd1 : 
                                        (_stream_conv2d_24_stream_oready && _stream_conv2d_24_sink_50_sink_wenable && (_stream_conv2d_24_sink_50_sink_sel == 21) && (write_rtl_bank_766 == 1))? 1'd1 : 0;
  assign ram_w8_l2048_id1_1_0_enable = (_stream_matmul_55_stream_oready && _stream_matmul_55_sink_26_sink_wenable && (_stream_matmul_55_sink_26_sink_sel == 5) && (write_rtl_bank_1811 == 1))? 1'd1 : 
                                       (_stream_conv2d_24_stream_oready && _stream_conv2d_24_sink_50_sink_wenable && (_stream_conv2d_24_sink_50_sink_sel == 21) && (write_rtl_bank_766 == 1))? 1'd1 : 0;
  assign ram_w8_l2048_id1_2_0_addr = (_stream_matmul_55_stream_oready && _stream_matmul_55_sink_26_sink_wenable && (_stream_matmul_55_sink_26_sink_sel == 5) && (write_rtl_bank_1811 == 2))? _stream_matmul_55_sink_26_sink_waddr >> 2 : 
                                     (_stream_conv2d_24_stream_oready && _stream_conv2d_24_sink_50_sink_wenable && (_stream_conv2d_24_sink_50_sink_sel == 21) && (write_rtl_bank_766 == 2))? _stream_conv2d_24_sink_50_sink_waddr >> 2 : 'hx;
  assign ram_w8_l2048_id1_2_0_wdata = (_stream_matmul_55_stream_oready && _stream_matmul_55_sink_26_sink_wenable && (_stream_matmul_55_sink_26_sink_sel == 5) && (write_rtl_bank_1811 == 2))? _stream_matmul_55_sink_26_sink_wdata : 
                                      (_stream_conv2d_24_stream_oready && _stream_conv2d_24_sink_50_sink_wenable && (_stream_conv2d_24_sink_50_sink_sel == 21) && (write_rtl_bank_766 == 2))? _stream_conv2d_24_sink_50_sink_wdata : 'hx;
  assign ram_w8_l2048_id1_2_0_wenable = (_stream_matmul_55_stream_oready && _stream_matmul_55_sink_26_sink_wenable && (_stream_matmul_55_sink_26_sink_sel == 5) && (write_rtl_bank_1811 == 2))? 1'd1 : 
                                        (_stream_conv2d_24_stream_oready && _stream_conv2d_24_sink_50_sink_wenable && (_stream_conv2d_24_sink_50_sink_sel == 21) && (write_rtl_bank_766 == 2))? 1'd1 : 0;
  assign ram_w8_l2048_id1_2_0_enable = (_stream_matmul_55_stream_oready && _stream_matmul_55_sink_26_sink_wenable && (_stream_matmul_55_sink_26_sink_sel == 5) && (write_rtl_bank_1811 == 2))? 1'd1 : 
                                       (_stream_conv2d_24_stream_oready && _stream_conv2d_24_sink_50_sink_wenable && (_stream_conv2d_24_sink_50_sink_sel == 21) && (write_rtl_bank_766 == 2))? 1'd1 : 0;
  assign ram_w8_l2048_id1_3_0_addr = (_stream_matmul_55_stream_oready && _stream_matmul_55_sink_26_sink_wenable && (_stream_matmul_55_sink_26_sink_sel == 5) && (write_rtl_bank_1811 == 3))? _stream_matmul_55_sink_26_sink_waddr >> 2 : 
                                     (_stream_conv2d_24_stream_oready && _stream_conv2d_24_sink_50_sink_wenable && (_stream_conv2d_24_sink_50_sink_sel == 21) && (write_rtl_bank_766 == 3))? _stream_conv2d_24_sink_50_sink_waddr >> 2 : 'hx;
  assign ram_w8_l2048_id1_3_0_wdata = (_stream_matmul_55_stream_oready && _stream_matmul_55_sink_26_sink_wenable && (_stream_matmul_55_sink_26_sink_sel == 5) && (write_rtl_bank_1811 == 3))? _stream_matmul_55_sink_26_sink_wdata : 
                                      (_stream_conv2d_24_stream_oready && _stream_conv2d_24_sink_50_sink_wenable && (_stream_conv2d_24_sink_50_sink_sel == 21) && (write_rtl_bank_766 == 3))? _stream_conv2d_24_sink_50_sink_wdata : 'hx;
  assign ram_w8_l2048_id1_3_0_wenable = (_stream_matmul_55_stream_oready && _stream_matmul_55_sink_26_sink_wenable && (_stream_matmul_55_sink_26_sink_sel == 5) && (write_rtl_bank_1811 == 3))? 1'd1 : 
                                        (_stream_conv2d_24_stream_oready && _stream_conv2d_24_sink_50_sink_wenable && (_stream_conv2d_24_sink_50_sink_sel == 21) && (write_rtl_bank_766 == 3))? 1'd1 : 0;
  assign ram_w8_l2048_id1_3_0_enable = (_stream_matmul_55_stream_oready && _stream_matmul_55_sink_26_sink_wenable && (_stream_matmul_55_sink_26_sink_sel == 5) && (write_rtl_bank_1811 == 3))? 1'd1 : 
                                       (_stream_conv2d_24_stream_oready && _stream_conv2d_24_sink_50_sink_wenable && (_stream_conv2d_24_sink_50_sink_sel == 21) && (write_rtl_bank_766 == 3))? 1'd1 : 0;
  reg [32-1:0] _stream_matmul_55_sink_26_sink_fsm_4;
  localparam _stream_matmul_55_sink_26_sink_fsm_4_init = 0;
  wire _set_flag_1812;
  assign _set_flag_1812 = matmul_55_comp_fsm == 4;
  assign _stream_matmul_55_run_flag = (_set_flag_1812)? 1 : 0;
  reg _tmp_1813;
  reg _tmp_1814;
  reg _tmp_1815;
  assign _add_tree_2_source_stop = _add_tree_2_stream_oready && 1'd0;
  reg _tmp_1816;
  reg _tmp_1817;
  assign _add_tree_2_sink_start = _tmp_1817;
  reg _tmp_1818;
  reg _tmp_1819;
  assign _add_tree_2_sink_stop = _tmp_1819;
  reg _tmp_1820;
  reg _tmp_1821;
  assign _add_tree_2_sink_busy = _tmp_1821;
  reg _tmp_1822;
  assign _add_tree_2_busy = _add_tree_2_source_busy || _add_tree_2_sink_busy || _add_tree_2_busy_reg;
  reg _tmp_1823;
  reg _tmp_1824;
  reg _tmp_1825;
  reg _tmp_1826;
  reg _tmp_1827;
  reg _tmp_1828;
  reg [1-1:0] __variable_wdata_941;
  assign stream_matmul_55__reduce_reset_data = __variable_wdata_941;
  reg _tmp_1829;
  reg _tmp_1830;
  reg _tmp_1831;
  reg _tmp_1832;
  assign _stream_matmul_55_source_stop = _stream_matmul_55_stream_oready && (_stream_matmul_55_source_11_idle && _stream_matmul_55_source_13_idle && _stream_matmul_55_source_15_idle && _stream_matmul_55_source_20_idle && _stream_matmul_55_source_21_idle && _stream_matmul_55_source_7_idle && _stream_matmul_55_source_9_idle && (_stream_matmul_55_fsm == 3));
  localparam _tmp_1833 = 1;
  wire [_tmp_1833-1:0] _tmp_1834;
  assign _tmp_1834 = _stream_matmul_55_source_11_idle && _stream_matmul_55_source_13_idle && _stream_matmul_55_source_15_idle && _stream_matmul_55_source_20_idle && _stream_matmul_55_source_21_idle && _stream_matmul_55_source_7_idle && _stream_matmul_55_source_9_idle && (_stream_matmul_55_fsm == 3);
  reg [_tmp_1833-1:0] _tmp_1835;
  localparam _tmp_1836 = 1;
  wire [_tmp_1836-1:0] _tmp_1837;
  assign _tmp_1837 = _stream_matmul_55_source_11_idle && _stream_matmul_55_source_13_idle && _stream_matmul_55_source_15_idle && _stream_matmul_55_source_20_idle && _stream_matmul_55_source_21_idle && _stream_matmul_55_source_7_idle && _stream_matmul_55_source_9_idle && (_stream_matmul_55_fsm == 3);
  reg [_tmp_1836-1:0] _tmp_1838;
  reg _tmp_1839;
  reg _tmp_1840;
  reg _tmp_1841;
  reg _tmp_1842;
  reg _tmp_1843;
  reg _tmp_1844;
  reg _tmp_1845;
  reg _tmp_1846;
  reg _tmp_1847;
  reg _tmp_1848;
  reg _tmp_1849;
  reg _tmp_1850;
  reg _tmp_1851;
  reg _tmp_1852;
  reg _tmp_1853;
  reg _tmp_1854;
  reg _tmp_1855;
  reg _tmp_1856;
  reg _tmp_1857;
  reg _tmp_1858;
  reg _tmp_1859;
  reg _tmp_1860;
  reg _tmp_1861;
  reg _tmp_1862;
  reg _tmp_1863;
  reg _tmp_1864;
  reg _tmp_1865;
  reg _tmp_1866;
  reg _tmp_1867;
  reg _tmp_1868;
  reg _tmp_1869;
  assign _stream_matmul_55_sink_start = _tmp_1869;
  reg _tmp_1870;
  reg _tmp_1871;
  reg _tmp_1872;
  reg _tmp_1873;
  reg _tmp_1874;
  reg _tmp_1875;
  reg _tmp_1876;
  reg _tmp_1877;
  reg _tmp_1878;
  reg _tmp_1879;
  reg _tmp_1880;
  reg _tmp_1881;
  reg _tmp_1882;
  reg _tmp_1883;
  reg _tmp_1884;
  reg _tmp_1885;
  reg _tmp_1886;
  reg _tmp_1887;
  reg _tmp_1888;
  reg _tmp_1889;
  reg _tmp_1890;
  reg _tmp_1891;
  reg _tmp_1892;
  reg _tmp_1893;
  reg _tmp_1894;
  reg _tmp_1895;
  reg _tmp_1896;
  reg _tmp_1897;
  reg _tmp_1898;
  reg _tmp_1899;
  reg _tmp_1900;
  assign _stream_matmul_55_sink_stop = _tmp_1900;
  reg _tmp_1901;
  reg _tmp_1902;
  reg _tmp_1903;
  reg _tmp_1904;
  reg _tmp_1905;
  reg _tmp_1906;
  reg _tmp_1907;
  reg _tmp_1908;
  reg _tmp_1909;
  reg _tmp_1910;
  reg _tmp_1911;
  reg _tmp_1912;
  reg _tmp_1913;
  reg _tmp_1914;
  reg _tmp_1915;
  reg _tmp_1916;
  reg _tmp_1917;
  reg _tmp_1918;
  reg _tmp_1919;
  reg _tmp_1920;
  reg _tmp_1921;
  reg _tmp_1922;
  reg _tmp_1923;
  reg _tmp_1924;
  reg _tmp_1925;
  reg _tmp_1926;
  reg _tmp_1927;
  reg _tmp_1928;
  reg _tmp_1929;
  reg _tmp_1930;
  reg _tmp_1931;
  assign _stream_matmul_55_sink_busy = _tmp_1931;
  reg _tmp_1932;
  assign _stream_matmul_55_busy = _stream_matmul_55_source_busy || _stream_matmul_55_sink_busy || _stream_matmul_55_busy_reg;
  wire matmul_55_dma_out_mask_0;
  assign matmul_55_dma_out_mask_0 = matmul_55_out_row_count + 0 >= cparam_matmul_55_out_num_row;
  wire [32-1:0] _dma_write_packed_high_local_size_1933;
  assign _dma_write_packed_high_local_size_1933 = matmul_55_next_out_write_size >> 2;
  wire [2-1:0] _dma_write_packed_low_local_size_1934;
  assign _dma_write_packed_low_local_size_1934 = matmul_55_next_out_write_size & { 2{ 1'd1 } };
  wire [32-1:0] _dma_write_packed_local_packed_size_1935;
  assign _dma_write_packed_local_packed_size_1935 = (_dma_write_packed_low_local_size_1934 > 0)? _dma_write_packed_high_local_size_1933 + 1 : _dma_write_packed_high_local_size_1933;
  wire [32-1:0] mask_addr_shifted_1936;
  assign mask_addr_shifted_1936 = matmul_55_objaddr + (matmul_55_out_base_offset + cparam_matmul_55_out_offset_values_0) + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_1937;
  assign mask_addr_masked_1937 = mask_addr_shifted_1936 << 2;
  wire matmul_55_update_filter;
  assign matmul_55_update_filter = (cparam_matmul_55_data_stationary == 0) && (matmul_55_row_count >= cparam_matmul_55_max_row_count) && (matmul_55_bat_count >= cparam_matmul_55_max_bat_count) || (cparam_matmul_55_data_stationary == 1) && !cparam_matmul_55_keep_filter;
  wire matmul_55_update_act;
  assign matmul_55_update_act = (cparam_matmul_55_data_stationary == 1) && (matmul_55_och_count >= cparam_matmul_55_max_och_count) || (cparam_matmul_55_data_stationary == 0);
  wire matmul_55_mux_next_dma_flag_0;
  assign matmul_55_mux_next_dma_flag_0 = (matmul_55_row_select == 0)? (matmul_55_row_count >= cparam_matmul_55_max_row_count)? 1 : cparam_matmul_55_dma_flag_conds_0 : 1'd0;

  always @(posedge CLK) begin
    _RESETN_inv_1 <= RESETN_inv;
    _RESETN_inv_2 <= _RESETN_inv_1;
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      maxi_awaddr <= 0;
      maxi_awlen <= 0;
      maxi_awvalid <= 0;
      _maxi_waddr_cond_0_1 <= 0;
    end else begin
      if(_maxi_waddr_cond_0_1) begin
        maxi_awvalid <= 0;
      end 
      if((_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (_maxi_outstanding_wcount < 6) && ((_maxi_outstanding_wcount < 6) && (maxi_awready || !maxi_awvalid))) begin
        maxi_awaddr <= _maxi_write_global_addr;
        maxi_awlen <= _maxi_write_cur_global_size - 1;
        maxi_awvalid <= 1;
      end 
      if((_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (_maxi_outstanding_wcount < 6) && ((_maxi_outstanding_wcount < 6) && (maxi_awready || !maxi_awvalid)) && (_maxi_write_cur_global_size == 0)) begin
        maxi_awvalid <= 0;
      end 
      _maxi_waddr_cond_0_1 <= 1;
      if(maxi_awvalid && !maxi_awready) begin
        maxi_awvalid <= maxi_awvalid;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      _maxi_wdata_sb_0 <= 0;
      _maxi_wvalid_sb_0 <= 0;
      _maxi_wlast_sb_0 <= 0;
      _maxi_wstrb_sb_0 <= 0;
      _maxi_wdata_cond_0_1 <= 0;
      _maxi_wdata_cond_1_1 <= 0;
      _maxi_wdata_cond_2_1 <= 0;
    end else begin
      if(_maxi_wdata_cond_0_1) begin
        _maxi_wvalid_sb_0 <= 0;
        _maxi_wlast_sb_0 <= 0;
      end 
      if(_maxi_wdata_cond_1_1) begin
        _maxi_wvalid_sb_0 <= 0;
        _maxi_wlast_sb_0 <= 0;
      end 
      if(_maxi_wdata_cond_2_1) begin
        _maxi_wvalid_sb_0 <= 0;
        _maxi_wlast_sb_0 <= 0;
      end 
      if((_maxi_write_op_sel_buf == 1) && read_burst_packed_rvalid_1308 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)) && (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0)) begin
        _maxi_wdata_sb_0 <= read_burst_packed_rdata_1326;
        _maxi_wvalid_sb_0 <= 1;
        _maxi_wlast_sb_0 <= read_burst_packed_rlast_1309 || (_maxi_write_size_buf == 1);
        _maxi_wstrb_sb_0 <= { 4{ 1'd1 } };
      end 
      _maxi_wdata_cond_0_1 <= 1;
      if(_maxi_wvalid_sb_0 && !_maxi_wready_sb_0) begin
        _maxi_wvalid_sb_0 <= _maxi_wvalid_sb_0;
        _maxi_wlast_sb_0 <= _maxi_wlast_sb_0;
      end 
      if((_maxi_write_op_sel_buf == 2) && read_burst_packed_rvalid_1456 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)) && (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0)) begin
        _maxi_wdata_sb_0 <= read_burst_packed_rdata_1474;
        _maxi_wvalid_sb_0 <= 1;
        _maxi_wlast_sb_0 <= read_burst_packed_rlast_1457 || (_maxi_write_size_buf == 1);
        _maxi_wstrb_sb_0 <= { 4{ 1'd1 } };
      end 
      _maxi_wdata_cond_1_1 <= 1;
      if(_maxi_wvalid_sb_0 && !_maxi_wready_sb_0) begin
        _maxi_wvalid_sb_0 <= _maxi_wvalid_sb_0;
        _maxi_wlast_sb_0 <= _maxi_wlast_sb_0;
      end 
      if((_maxi_write_op_sel_buf == 3) && read_burst_packed_rvalid_1608 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)) && (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0)) begin
        _maxi_wdata_sb_0 <= read_burst_packed_rdata_1626;
        _maxi_wvalid_sb_0 <= 1;
        _maxi_wlast_sb_0 <= read_burst_packed_rlast_1609 || (_maxi_write_size_buf == 1);
        _maxi_wstrb_sb_0 <= { 4{ 1'd1 } };
      end 
      _maxi_wdata_cond_2_1 <= 1;
      if(_maxi_wvalid_sb_0 && !_maxi_wready_sb_0) begin
        _maxi_wvalid_sb_0 <= _maxi_wvalid_sb_0;
        _maxi_wlast_sb_0 <= _maxi_wlast_sb_0;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      _sb_maxi_writedata_data_6 <= 0;
      _sb_maxi_writedata_valid_7 <= 0;
      _sb_maxi_writedata_tmp_data_9 <= 0;
      _sb_maxi_writedata_tmp_valid_10 <= 0;
    end else begin
      if(_sb_maxi_writedata_m_ready_5 || !_sb_maxi_writedata_valid_7) begin
        _sb_maxi_writedata_data_6 <= _sb_maxi_writedata_next_data_11;
        _sb_maxi_writedata_valid_7 <= _sb_maxi_writedata_next_valid_12;
      end 
      if(!_sb_maxi_writedata_tmp_valid_10 && _sb_maxi_writedata_valid_7 && !_sb_maxi_writedata_m_ready_5) begin
        _sb_maxi_writedata_tmp_data_9 <= _sb_maxi_writedata_s_data_3;
        _sb_maxi_writedata_tmp_valid_10 <= _sb_maxi_writedata_s_valid_4;
      end 
      if(_sb_maxi_writedata_tmp_valid_10 && _sb_maxi_writedata_m_ready_5) begin
        _sb_maxi_writedata_tmp_valid_10 <= 0;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      maxi_araddr <= 0;
      maxi_arlen <= 0;
      maxi_arvalid <= 0;
      _maxi_raddr_cond_0_1 <= 0;
    end else begin
      if(_maxi_raddr_cond_0_1) begin
        maxi_arvalid <= 0;
      end 
      if((_maxi_read_req_fsm == 1) && (maxi_arready || !maxi_arvalid)) begin
        maxi_araddr <= _maxi_read_global_addr;
        maxi_arlen <= _maxi_read_cur_global_size - 1;
        maxi_arvalid <= 1;
      end 
      _maxi_raddr_cond_0_1 <= 1;
      if(maxi_arvalid && !maxi_arready) begin
        maxi_arvalid <= maxi_arvalid;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      _sb_maxi_readdata_data_21 <= 0;
      _sb_maxi_readdata_valid_22 <= 0;
      _sb_maxi_readdata_tmp_data_24 <= 0;
      _sb_maxi_readdata_tmp_valid_25 <= 0;
    end else begin
      if(_sb_maxi_readdata_m_ready_20 || !_sb_maxi_readdata_valid_22) begin
        _sb_maxi_readdata_data_21 <= _sb_maxi_readdata_next_data_26;
        _sb_maxi_readdata_valid_22 <= _sb_maxi_readdata_next_valid_27;
      end 
      if(!_sb_maxi_readdata_tmp_valid_25 && _sb_maxi_readdata_valid_22 && !_sb_maxi_readdata_m_ready_20) begin
        _sb_maxi_readdata_tmp_data_24 <= _sb_maxi_readdata_s_data_18;
        _sb_maxi_readdata_tmp_valid_25 <= _sb_maxi_readdata_s_valid_19;
      end 
      if(_sb_maxi_readdata_tmp_valid_25 && _sb_maxi_readdata_m_ready_20) begin
        _sb_maxi_readdata_tmp_valid_25 <= 0;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      _maxi_outstanding_wcount <= 0;
      _maxi_read_start <= 0;
      _maxi_write_start <= 0;
      _maxi_global_base_addr <= 0;
      _maxi_read_op_sel <= 0;
      _maxi_read_global_addr <= 0;
      _maxi_read_global_size <= 0;
      _maxi_read_local_addr <= 0;
      _maxi_read_local_stride <= 0;
      _maxi_read_local_size <= 0;
      _maxi_read_local_blocksize <= 0;
      _maxi_read_req_busy <= 0;
      _maxi_read_cur_global_size <= 0;
      _maxi_read_data_busy <= 0;
      _maxi_read_op_sel_buf <= 0;
      _maxi_read_local_addr_buf <= 0;
      _maxi_read_local_stride_buf <= 0;
      _maxi_read_local_size_buf <= 0;
      _maxi_read_local_blocksize_buf <= 0;
      _maxi_write_op_sel <= 0;
      _maxi_write_global_addr <= 0;
      _maxi_write_global_size <= 0;
      _maxi_write_local_addr <= 0;
      _maxi_write_local_stride <= 0;
      _maxi_write_local_size <= 0;
      _maxi_write_local_blocksize <= 0;
      _maxi_write_req_busy <= 0;
      _maxi_write_cur_global_size <= 0;
      _maxi_write_data_busy <= 0;
      _maxi_write_op_sel_buf <= 0;
      _maxi_write_local_addr_buf <= 0;
      _maxi_write_local_stride_buf <= 0;
      _maxi_write_size_buf <= 0;
      _maxi_write_local_blocksize_buf <= 0;
    end else begin
      if(maxi_awvalid && maxi_awready && !(maxi_bvalid && maxi_bready) && (_maxi_outstanding_wcount < 7)) begin
        _maxi_outstanding_wcount <= _maxi_outstanding_wcount + 1;
      end 
      if(!(maxi_awvalid && maxi_awready) && (maxi_bvalid && maxi_bready) && (_maxi_outstanding_wcount > 0)) begin
        _maxi_outstanding_wcount <= _maxi_outstanding_wcount - 1;
      end 
      _maxi_read_start <= 0;
      _maxi_write_start <= 0;
      _maxi_global_base_addr <= _saxi_register_32;
      if((control_conv2d_24 == 2) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 1;
        _maxi_read_global_addr <= mask_addr_masked_55;
        _maxi_read_global_size <= cparam_conv2d_24_bias_num;
        _maxi_read_local_addr <= 0;
        _maxi_read_local_stride <= 1;
        _maxi_read_local_size <= cparam_conv2d_24_bias_num;
        _maxi_read_local_blocksize <= 1;
      end 
      if((_maxi_read_req_fsm == 0) && _maxi_read_start) begin
        _maxi_read_req_busy <= 1;
      end 
      if(_maxi_read_start && _maxi_read_req_fifo_almost_full) begin
        _maxi_read_start <= 1;
      end 
      if((_maxi_read_req_fsm == 0) && (_maxi_read_start || _maxi_read_cont) && !_maxi_read_req_fifo_almost_full && (_maxi_read_global_size <= 256) && ((mask_addr_masked_65 & 4095) + (_maxi_read_global_size << 2) >= 4096)) begin
        _maxi_read_cur_global_size <= 4096 - (mask_addr_masked_67 & 4095) >> 2;
        _maxi_read_global_size <= _maxi_read_global_size - (4096 - (mask_addr_masked_69 & 4095) >> 2);
      end else if((_maxi_read_req_fsm == 0) && (_maxi_read_start || _maxi_read_cont) && !_maxi_read_req_fifo_almost_full && (_maxi_read_global_size <= 256)) begin
        _maxi_read_cur_global_size <= _maxi_read_global_size;
        _maxi_read_global_size <= 0;
      end else if((_maxi_read_req_fsm == 0) && (_maxi_read_start || _maxi_read_cont) && !_maxi_read_req_fifo_almost_full && ((mask_addr_masked_71 & 4095) + 1024 >= 4096)) begin
        _maxi_read_cur_global_size <= 4096 - (mask_addr_masked_73 & 4095) >> 2;
        _maxi_read_global_size <= _maxi_read_global_size - (4096 - (mask_addr_masked_75 & 4095) >> 2);
      end else if((_maxi_read_req_fsm == 0) && (_maxi_read_start || _maxi_read_cont) && !_maxi_read_req_fifo_almost_full) begin
        _maxi_read_cur_global_size <= 256;
        _maxi_read_global_size <= _maxi_read_global_size - 256;
      end 
      if((_maxi_read_req_fsm == 1) && (maxi_arready || !maxi_arvalid)) begin
        _maxi_read_global_addr <= _maxi_read_global_addr + (_maxi_read_cur_global_size << 2);
      end 
      if((_maxi_read_req_fsm == 1) && (maxi_arready || !maxi_arvalid) && (_maxi_read_global_size == 0)) begin
        _maxi_read_req_busy <= 0;
      end 
      if((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 1))) begin
        _maxi_read_data_busy <= 1;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_busy <= 0;
      end 
      if((control_conv2d_24 == 4) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 2;
        _maxi_read_global_addr <= mask_addr_masked_84;
        _maxi_read_global_size <= _dma_read_packed_local_packed_size_82;
        _maxi_read_local_addr <= 0;
        _maxi_read_local_stride <= 4;
        _maxi_read_local_size <= _dma_read_packed_local_packed_size_82;
        _maxi_read_local_blocksize <= 1;
      end 
      if((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 2))) begin
        _maxi_read_data_busy <= 1;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_busy <= 0;
      end 
      if((control_conv2d_24 == 8) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 3;
        _maxi_read_global_addr <= mask_addr_masked_104;
        _maxi_read_global_size <= _dma_write_block_local_size_99;
        _maxi_read_local_addr <= conv2d_24_filter_page_dma_offset;
        _maxi_read_local_stride <= 4;
        _maxi_read_local_size <= _dma_write_block_local_size_99;
        _maxi_read_local_blocksize <= _dma_read_block_local_blocksize_102;
      end 
      if((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 3))) begin
        _maxi_read_data_busy <= 1;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_busy <= 0;
      end 
      if((control_conv2d_24 == 14) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 4;
        _maxi_read_global_addr <= mask_addr_masked_242;
        _maxi_read_global_size <= _dma_write_block_local_size_237;
        _maxi_read_local_addr <= conv2d_24_act_page_dma_offset_0;
        _maxi_read_local_stride <= 4;
        _maxi_read_local_size <= _dma_write_block_local_size_237;
        _maxi_read_local_blocksize <= _dma_read_block_local_blocksize_240;
      end 
      if((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 4))) begin
        _maxi_read_data_busy <= 1;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_busy <= 0;
      end 
      if((control_conv2d_24 == 17) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 5;
        _maxi_read_global_addr <= mask_addr_masked_296;
        _maxi_read_global_size <= _dma_write_block_local_size_291;
        _maxi_read_local_addr <= conv2d_24_act_page_dma_offset_1;
        _maxi_read_local_stride <= 4;
        _maxi_read_local_size <= _dma_write_block_local_size_291;
        _maxi_read_local_blocksize <= _dma_read_block_local_blocksize_294;
      end 
      if((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 5))) begin
        _maxi_read_data_busy <= 1;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_busy <= 0;
      end 
      if((control_conv2d_24 == 20) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 6;
        _maxi_read_global_addr <= mask_addr_masked_350;
        _maxi_read_global_size <= _dma_write_block_local_size_345;
        _maxi_read_local_addr <= conv2d_24_act_page_dma_offset_2;
        _maxi_read_local_stride <= 4;
        _maxi_read_local_size <= _dma_write_block_local_size_345;
        _maxi_read_local_blocksize <= _dma_read_block_local_blocksize_348;
      end 
      if((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 6))) begin
        _maxi_read_data_busy <= 1;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_busy <= 0;
      end 
      if((control_conv2d_24 == 29) && _maxi_write_req_idle) begin
        _maxi_write_start <= 1;
        _maxi_write_op_sel <= 1;
        _maxi_write_global_addr <= mask_addr_masked_1276;
        _maxi_write_global_size <= _dma_write_packed_local_packed_size_1274;
        _maxi_write_local_addr <= conv2d_24_out_laddr_offset + conv2d_24_out_page_dma_offset;
        _maxi_write_local_stride <= 4;
        _maxi_write_local_size <= _dma_write_packed_local_packed_size_1274;
        _maxi_write_local_blocksize <= 1;
      end 
      if((_maxi_write_req_fsm == 0) && _maxi_write_start) begin
        _maxi_write_req_busy <= 1;
      end 
      if(_maxi_write_start && _maxi_write_req_fifo_almost_full) begin
        _maxi_write_start <= 1;
      end 
      if((_maxi_write_req_fsm == 0) && (_maxi_write_start || _maxi_write_cont) && !_maxi_write_req_fifo_almost_full && (_maxi_write_global_size <= 256) && ((mask_addr_masked_1286 & 4095) + (_maxi_write_global_size << 2) >= 4096)) begin
        _maxi_write_cur_global_size <= 4096 - (mask_addr_masked_1288 & 4095) >> 2;
        _maxi_write_global_size <= _maxi_write_global_size - (4096 - (mask_addr_masked_1290 & 4095) >> 2);
      end else if((_maxi_write_req_fsm == 0) && (_maxi_write_start || _maxi_write_cont) && !_maxi_write_req_fifo_almost_full && (_maxi_write_global_size <= 256)) begin
        _maxi_write_cur_global_size <= _maxi_write_global_size;
        _maxi_write_global_size <= 0;
      end else if((_maxi_write_req_fsm == 0) && (_maxi_write_start || _maxi_write_cont) && !_maxi_write_req_fifo_almost_full && ((mask_addr_masked_1292 & 4095) + 1024 >= 4096)) begin
        _maxi_write_cur_global_size <= 4096 - (mask_addr_masked_1294 & 4095) >> 2;
        _maxi_write_global_size <= _maxi_write_global_size - (4096 - (mask_addr_masked_1296 & 4095) >> 2);
      end else if((_maxi_write_req_fsm == 0) && (_maxi_write_start || _maxi_write_cont) && !_maxi_write_req_fifo_almost_full) begin
        _maxi_write_cur_global_size <= 256;
        _maxi_write_global_size <= _maxi_write_global_size - 256;
      end 
      if((_maxi_write_req_fsm == 1) && ((_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (maxi_awready || !maxi_awvalid) && (_maxi_outstanding_wcount < 6))) begin
        _maxi_write_global_addr <= _maxi_write_global_addr + (_maxi_write_cur_global_size << 2);
      end 
      if((_maxi_write_req_fsm == 1) && ((_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (maxi_awready || !maxi_awvalid) && (_maxi_outstanding_wcount < 6)) && (_maxi_write_global_size == 0)) begin
        _maxi_write_req_busy <= 0;
      end 
      if((_maxi_write_data_fsm == 0) && (!_maxi_write_data_busy && !_maxi_write_req_fifo_empty && (_maxi_write_op_sel_fifo == 1))) begin
        _maxi_write_data_busy <= 1;
        _maxi_write_op_sel_buf <= _maxi_write_op_sel_fifo;
        _maxi_write_local_addr_buf <= _maxi_write_local_addr_fifo;
        _maxi_write_local_stride_buf <= _maxi_write_local_stride_fifo;
        _maxi_write_size_buf <= _maxi_write_size_fifo;
        _maxi_write_local_blocksize_buf <= _maxi_write_local_blocksize_fifo;
      end 
      if(_maxi_write_data_fsm == 1) begin
        _maxi_write_size_buf <= 0;
      end 
      if((_maxi_write_data_fsm == 2) && (!_maxi_write_req_fifo_empty && (_maxi_write_size_buf == 0))) begin
        _maxi_write_size_buf <= _maxi_write_size_fifo;
      end 
      if((_maxi_write_data_fsm == 2) && read_burst_packed_rvalid_1308 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) begin
        _maxi_write_size_buf <= _maxi_write_size_buf - 1;
      end 
      if((_maxi_write_data_fsm == 2) && ((_maxi_write_op_sel_buf == 1) && read_burst_packed_rvalid_1308 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) && read_burst_packed_rlast_1309) begin
        _maxi_write_data_busy <= 0;
      end 
      if((control_max_pool_serial_26 == 5) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 7;
        _maxi_read_global_addr <= mask_addr_masked_1331;
        _maxi_read_global_size <= _dma_read_packed_local_packed_size_1329;
        _maxi_read_local_addr <= max_pool_serial_26_act_page_dma_offset;
        _maxi_read_local_stride <= 4;
        _maxi_read_local_size <= _dma_read_packed_local_packed_size_1329;
        _maxi_read_local_blocksize <= 1;
      end 
      if((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 7))) begin
        _maxi_read_data_busy <= 1;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_busy <= 0;
      end 
      if((control_max_pool_serial_26 == 8) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 7;
        _maxi_read_global_addr <= mask_addr_masked_1348;
        _maxi_read_global_size <= _dma_read_packed_local_packed_size_1346;
        _maxi_read_local_addr <= max_pool_serial_26_act_page_dma_offset + cparam_max_pool_serial_26_act_read_size;
        _maxi_read_local_stride <= 4;
        _maxi_read_local_size <= _dma_read_packed_local_packed_size_1346;
        _maxi_read_local_blocksize <= 1;
      end 
      if((control_max_pool_serial_26 == 15) && _maxi_write_req_idle) begin
        _maxi_write_start <= 1;
        _maxi_write_op_sel <= 2;
        _maxi_write_global_addr <= mask_addr_masked_1452;
        _maxi_write_global_size <= _dma_write_packed_local_packed_size_1450;
        _maxi_write_local_addr <= max_pool_serial_26_out_page_dma_offset;
        _maxi_write_local_stride <= 4;
        _maxi_write_local_size <= _dma_write_packed_local_packed_size_1450;
        _maxi_write_local_blocksize <= 1;
      end 
      if((_maxi_write_data_fsm == 0) && (!_maxi_write_data_busy && !_maxi_write_req_fifo_empty && (_maxi_write_op_sel_fifo == 2))) begin
        _maxi_write_data_busy <= 1;
        _maxi_write_op_sel_buf <= _maxi_write_op_sel_fifo;
        _maxi_write_local_addr_buf <= _maxi_write_local_addr_fifo;
        _maxi_write_local_stride_buf <= _maxi_write_local_stride_fifo;
        _maxi_write_size_buf <= _maxi_write_size_fifo;
        _maxi_write_local_blocksize_buf <= _maxi_write_local_blocksize_fifo;
      end 
      if(_maxi_write_data_fsm == 1) begin
        _maxi_write_size_buf <= 0;
      end 
      if((_maxi_write_data_fsm == 2) && (!_maxi_write_req_fifo_empty && (_maxi_write_size_buf == 0))) begin
        _maxi_write_size_buf <= _maxi_write_size_fifo;
      end 
      if((_maxi_write_data_fsm == 2) && read_burst_packed_rvalid_1456 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) begin
        _maxi_write_size_buf <= _maxi_write_size_buf - 1;
      end 
      if((_maxi_write_data_fsm == 2) && ((_maxi_write_op_sel_buf == 2) && read_burst_packed_rvalid_1456 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) && read_burst_packed_rlast_1457) begin
        _maxi_write_data_busy <= 0;
      end 
      if((control_avg_pool_serial_52 == 5) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 8;
        _maxi_read_global_addr <= mask_addr_masked_1479;
        _maxi_read_global_size <= _dma_read_packed_local_packed_size_1477;
        _maxi_read_local_addr <= avg_pool_serial_52_act_page_dma_offset;
        _maxi_read_local_stride <= 4;
        _maxi_read_local_size <= _dma_read_packed_local_packed_size_1477;
        _maxi_read_local_blocksize <= 1;
      end 
      if((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 8))) begin
        _maxi_read_data_busy <= 1;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_busy <= 0;
      end 
      if((control_avg_pool_serial_52 == 12) && _maxi_write_req_idle) begin
        _maxi_write_start <= 1;
        _maxi_write_op_sel <= 3;
        _maxi_write_global_addr <= mask_addr_masked_1604;
        _maxi_write_global_size <= _dma_write_packed_local_packed_size_1602;
        _maxi_write_local_addr <= avg_pool_serial_52_out_page_dma_offset;
        _maxi_write_local_stride <= 4;
        _maxi_write_local_size <= _dma_write_packed_local_packed_size_1602;
        _maxi_write_local_blocksize <= 1;
      end 
      if((_maxi_write_data_fsm == 0) && (!_maxi_write_data_busy && !_maxi_write_req_fifo_empty && (_maxi_write_op_sel_fifo == 3))) begin
        _maxi_write_data_busy <= 1;
        _maxi_write_op_sel_buf <= _maxi_write_op_sel_fifo;
        _maxi_write_local_addr_buf <= _maxi_write_local_addr_fifo;
        _maxi_write_local_stride_buf <= _maxi_write_local_stride_fifo;
        _maxi_write_size_buf <= _maxi_write_size_fifo;
        _maxi_write_local_blocksize_buf <= _maxi_write_local_blocksize_fifo;
      end 
      if(_maxi_write_data_fsm == 1) begin
        _maxi_write_size_buf <= 0;
      end 
      if((_maxi_write_data_fsm == 2) && (!_maxi_write_req_fifo_empty && (_maxi_write_size_buf == 0))) begin
        _maxi_write_size_buf <= _maxi_write_size_fifo;
      end 
      if((_maxi_write_data_fsm == 2) && read_burst_packed_rvalid_1608 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) begin
        _maxi_write_size_buf <= _maxi_write_size_buf - 1;
      end 
      if((_maxi_write_data_fsm == 2) && ((_maxi_write_op_sel_buf == 3) && read_burst_packed_rvalid_1608 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) && read_burst_packed_rlast_1609) begin
        _maxi_write_data_busy <= 0;
      end 
      if((control_matmul_55 == 2) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 1;
        _maxi_read_global_addr <= mask_addr_masked_1628;
        _maxi_read_global_size <= cparam_matmul_55_bias_num;
        _maxi_read_local_addr <= 0;
        _maxi_read_local_stride <= 1;
        _maxi_read_local_size <= cparam_matmul_55_bias_num;
        _maxi_read_local_blocksize <= 1;
      end 
      if((control_matmul_55 == 4) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 2;
        _maxi_read_global_addr <= mask_addr_masked_1633;
        _maxi_read_global_size <= _dma_read_packed_local_packed_size_1631;
        _maxi_read_local_addr <= 0;
        _maxi_read_local_stride <= 4;
        _maxi_read_local_size <= _dma_read_packed_local_packed_size_1631;
        _maxi_read_local_blocksize <= 1;
      end 
      if((control_matmul_55 == 8) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 7;
        _maxi_read_global_addr <= mask_addr_masked_1638;
        _maxi_read_global_size <= _dma_read_packed_local_packed_size_1636;
        _maxi_read_local_addr <= matmul_55_filter_page_dma_offset;
        _maxi_read_local_stride <= 4;
        _maxi_read_local_size <= _dma_read_packed_local_packed_size_1636;
        _maxi_read_local_blocksize <= 1;
      end 
      if((control_matmul_55 == 14) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 9;
        _maxi_read_global_addr <= mask_addr_masked_1643;
        _maxi_read_global_size <= _dma_read_packed_local_packed_size_1641;
        _maxi_read_local_addr <= matmul_55_act_page_dma_offset_0;
        _maxi_read_local_stride <= 4;
        _maxi_read_local_size <= _dma_read_packed_local_packed_size_1641;
        _maxi_read_local_blocksize <= 1;
      end 
      if((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 9))) begin
        _maxi_read_data_busy <= 1;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_busy <= 0;
      end 
      if((control_matmul_55 == 23) && _maxi_write_req_idle) begin
        _maxi_write_start <= 1;
        _maxi_write_op_sel <= 1;
        _maxi_write_global_addr <= mask_addr_masked_1937;
        _maxi_write_global_size <= _dma_write_packed_local_packed_size_1935;
        _maxi_write_local_addr <= matmul_55_out_laddr_offset + matmul_55_out_page_dma_offset;
        _maxi_write_local_stride <= 4;
        _maxi_write_local_size <= _dma_write_packed_local_packed_size_1935;
        _maxi_write_local_blocksize <= 1;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      count__maxi_read_req_fifo <= 0;
      __tmp_63_1 <= 0;
    end else begin
      if(_maxi_read_req_fifo_enq && !_maxi_read_req_fifo_full && (_maxi_read_req_fifo_deq && !_maxi_read_req_fifo_empty)) begin
        count__maxi_read_req_fifo <= count__maxi_read_req_fifo;
      end else if(_maxi_read_req_fifo_enq && !_maxi_read_req_fifo_full) begin
        count__maxi_read_req_fifo <= count__maxi_read_req_fifo + 1;
      end else if(_maxi_read_req_fifo_deq && !_maxi_read_req_fifo_empty) begin
        count__maxi_read_req_fifo <= count__maxi_read_req_fifo - 1;
      end 
      __tmp_63_1 <= _tmp_63;
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      count__maxi_write_req_fifo <= 0;
      __tmp_1284_1 <= 0;
      __tmp_1304_1 <= 0;
    end else begin
      if(_maxi_write_req_fifo_enq && !_maxi_write_req_fifo_full && (_maxi_write_req_fifo_deq && !_maxi_write_req_fifo_empty)) begin
        count__maxi_write_req_fifo <= count__maxi_write_req_fifo;
      end else if(_maxi_write_req_fifo_enq && !_maxi_write_req_fifo_full) begin
        count__maxi_write_req_fifo <= count__maxi_write_req_fifo + 1;
      end else if(_maxi_write_req_fifo_deq && !_maxi_write_req_fifo_empty) begin
        count__maxi_write_req_fifo <= count__maxi_write_req_fifo - 1;
      end 
      __tmp_1284_1 <= _tmp_1284;
      __tmp_1304_1 <= _tmp_1304;
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      saxi_rdata <= 0;
      saxi_rvalid <= 0;
      _saxi_rdata_cond_0_1 <= 0;
    end else begin
      if(_saxi_rdata_cond_0_1) begin
        saxi_rvalid <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid)) begin
        saxi_rdata <= axislite_rdata_46;
        saxi_rvalid <= 1;
      end 
      _saxi_rdata_cond_0_1 <= 1;
      if(saxi_rvalid && !saxi_rready) begin
        saxi_rvalid <= saxi_rvalid;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      saxi_bvalid <= 0;
      prev_awvalid_43 <= 0;
      prev_arvalid_44 <= 0;
      writevalid_41 <= 0;
      readvalid_42 <= 0;
      addr_40 <= 0;
      _saxi_register_0 <= 0;
      _saxi_flag_0 <= 0;
      _saxi_register_1 <= 0;
      _saxi_flag_1 <= 0;
      _saxi_register_2 <= 0;
      _saxi_flag_2 <= 0;
      _saxi_register_3 <= 0;
      _saxi_flag_3 <= 0;
      _saxi_register_4 <= 0;
      _saxi_flag_4 <= 0;
      _saxi_register_5 <= 0;
      _saxi_flag_5 <= 0;
      _saxi_register_6 <= 0;
      _saxi_flag_6 <= 0;
      _saxi_register_7 <= 0;
      _saxi_flag_7 <= 0;
      _saxi_register_8 <= 0;
      _saxi_flag_8 <= 0;
      _saxi_register_9 <= 0;
      _saxi_flag_9 <= 0;
      _saxi_register_10 <= 0;
      _saxi_flag_10 <= 0;
      _saxi_register_11 <= 0;
      _saxi_flag_11 <= 0;
      _saxi_register_12 <= 0;
      _saxi_flag_12 <= 0;
      _saxi_register_13 <= 0;
      _saxi_flag_13 <= 0;
      _saxi_register_14 <= 0;
      _saxi_flag_14 <= 0;
      _saxi_register_15 <= 0;
      _saxi_flag_15 <= 0;
      _saxi_register_16 <= 0;
      _saxi_flag_16 <= 0;
      _saxi_register_17 <= 0;
      _saxi_flag_17 <= 0;
      _saxi_register_18 <= 0;
      _saxi_flag_18 <= 0;
      _saxi_register_19 <= 0;
      _saxi_flag_19 <= 0;
      _saxi_register_20 <= 0;
      _saxi_flag_20 <= 0;
      _saxi_register_21 <= 0;
      _saxi_flag_21 <= 0;
      _saxi_register_22 <= 0;
      _saxi_flag_22 <= 0;
      _saxi_register_23 <= 0;
      _saxi_flag_23 <= 0;
      _saxi_register_24 <= 0;
      _saxi_flag_24 <= 0;
      _saxi_register_25 <= 0;
      _saxi_flag_25 <= 0;
      _saxi_register_26 <= 0;
      _saxi_flag_26 <= 0;
      _saxi_register_27 <= 0;
      _saxi_flag_27 <= 0;
      _saxi_register_28 <= 0;
      _saxi_flag_28 <= 0;
      _saxi_register_29 <= 0;
      _saxi_flag_29 <= 0;
      _saxi_register_30 <= 0;
      _saxi_flag_30 <= 0;
      _saxi_register_31 <= 142091904;
      _saxi_flag_31 <= 0;
      _saxi_register_32 <= 0;
      _saxi_flag_32 <= 0;
      _saxi_register_33 <= 133102208;
      _saxi_flag_33 <= 0;
      _saxi_register_34 <= 0;
      _saxi_flag_34 <= 0;
      _saxi_register_35 <= 1024;
      _saxi_flag_35 <= 0;
      _saxi_register_36 <= 201728;
      _saxi_flag_36 <= 0;
      _saxi_register_11[0] <= (0 >> 0) & 1'd1;
      _saxi_register_9[0] <= (0 >> 0) & 1'd1;
      _saxi_register_11[1] <= (0 >> 1) & 1'd1;
      _saxi_register_9[1] <= (0 >> 1) & 1'd1;
      _saxi_register_11[2] <= (0 >> 2) & 1'd1;
      _saxi_register_9[2] <= (0 >> 2) & 1'd1;
      _saxi_register_11[3] <= (0 >> 3) & 1'd1;
      _saxi_register_9[3] <= (0 >> 3) & 1'd1;
      _saxi_register_11[4] <= (0 >> 4) & 1'd1;
      _saxi_register_9[4] <= (0 >> 4) & 1'd1;
      _saxi_register_11[5] <= (0 >> 5) & 1'd1;
      _saxi_register_9[5] <= (0 >> 5) & 1'd1;
      _saxi_register_11[6] <= (0 >> 6) & 1'd1;
      _saxi_register_9[6] <= (0 >> 6) & 1'd1;
      _saxi_register_11[7] <= (0 >> 7) & 1'd1;
      _saxi_register_9[7] <= (0 >> 7) & 1'd1;
      _saxi_register_11[8] <= (0 >> 8) & 1'd1;
      _saxi_register_9[8] <= (0 >> 8) & 1'd1;
      _saxi_register_11[9] <= (0 >> 9) & 1'd1;
      _saxi_register_9[9] <= (0 >> 9) & 1'd1;
      _saxi_register_11[10] <= (0 >> 10) & 1'd1;
      _saxi_register_9[10] <= (0 >> 10) & 1'd1;
      _saxi_register_11[11] <= (0 >> 11) & 1'd1;
      _saxi_register_9[11] <= (0 >> 11) & 1'd1;
      _saxi_register_11[12] <= (0 >> 12) & 1'd1;
      _saxi_register_9[12] <= (0 >> 12) & 1'd1;
      _saxi_register_11[13] <= (0 >> 13) & 1'd1;
      _saxi_register_9[13] <= (0 >> 13) & 1'd1;
      _saxi_register_11[14] <= (0 >> 14) & 1'd1;
      _saxi_register_9[14] <= (0 >> 14) & 1'd1;
      _saxi_register_11[15] <= (0 >> 15) & 1'd1;
      _saxi_register_9[15] <= (0 >> 15) & 1'd1;
      _saxi_register_11[16] <= (0 >> 16) & 1'd1;
      _saxi_register_9[16] <= (0 >> 16) & 1'd1;
      _saxi_register_11[17] <= (0 >> 17) & 1'd1;
      _saxi_register_9[17] <= (0 >> 17) & 1'd1;
      _saxi_register_11[18] <= (0 >> 18) & 1'd1;
      _saxi_register_9[18] <= (0 >> 18) & 1'd1;
      _saxi_register_11[19] <= (0 >> 19) & 1'd1;
      _saxi_register_9[19] <= (0 >> 19) & 1'd1;
      _saxi_register_11[20] <= (0 >> 20) & 1'd1;
      _saxi_register_9[20] <= (0 >> 20) & 1'd1;
      _saxi_register_11[21] <= (0 >> 21) & 1'd1;
      _saxi_register_9[21] <= (0 >> 21) & 1'd1;
      _saxi_register_11[22] <= (0 >> 22) & 1'd1;
      _saxi_register_9[22] <= (0 >> 22) & 1'd1;
      _saxi_register_11[23] <= (0 >> 23) & 1'd1;
      _saxi_register_9[23] <= (0 >> 23) & 1'd1;
      _saxi_register_11[24] <= (0 >> 24) & 1'd1;
      _saxi_register_9[24] <= (0 >> 24) & 1'd1;
      _saxi_register_11[25] <= (0 >> 25) & 1'd1;
      _saxi_register_9[25] <= (0 >> 25) & 1'd1;
      _saxi_register_11[26] <= (0 >> 26) & 1'd1;
      _saxi_register_9[26] <= (0 >> 26) & 1'd1;
      _saxi_register_11[27] <= (0 >> 27) & 1'd1;
      _saxi_register_9[27] <= (0 >> 27) & 1'd1;
      _saxi_register_11[28] <= (0 >> 28) & 1'd1;
      _saxi_register_9[28] <= (0 >> 28) & 1'd1;
      _saxi_register_11[29] <= (0 >> 29) & 1'd1;
      _saxi_register_9[29] <= (0 >> 29) & 1'd1;
      _saxi_register_11[30] <= (0 >> 30) & 1'd1;
      _saxi_register_9[30] <= (0 >> 30) & 1'd1;
      _saxi_register_11[31] <= (0 >> 31) & 1'd1;
      _saxi_register_9[31] <= (0 >> 31) & 1'd1;
      internal_state_counter <= 0;
    end else begin
      if(saxi_bvalid && saxi_bready) begin
        saxi_bvalid <= 0;
      end 
      if(saxi_wvalid && saxi_wready) begin
        saxi_bvalid <= 1;
      end 
      prev_awvalid_43 <= saxi_awvalid;
      prev_arvalid_44 <= saxi_arvalid;
      writevalid_41 <= 0;
      readvalid_42 <= 0;
      if(saxi_awready && saxi_awvalid && !saxi_bvalid) begin
        addr_40 <= saxi_awaddr;
        writevalid_41 <= 1;
      end else if(saxi_arready && saxi_arvalid) begin
        addr_40 <= saxi_araddr;
        readvalid_42 <= 1;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 0)) begin
        _saxi_register_0 <= axislite_resetval_48;
        _saxi_flag_0 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 1)) begin
        _saxi_register_1 <= axislite_resetval_48;
        _saxi_flag_1 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 2)) begin
        _saxi_register_2 <= axislite_resetval_48;
        _saxi_flag_2 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 3)) begin
        _saxi_register_3 <= axislite_resetval_48;
        _saxi_flag_3 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 4)) begin
        _saxi_register_4 <= axislite_resetval_48;
        _saxi_flag_4 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 5)) begin
        _saxi_register_5 <= axislite_resetval_48;
        _saxi_flag_5 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 6)) begin
        _saxi_register_6 <= axislite_resetval_48;
        _saxi_flag_6 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 7)) begin
        _saxi_register_7 <= axislite_resetval_48;
        _saxi_flag_7 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 8)) begin
        _saxi_register_8 <= axislite_resetval_48;
        _saxi_flag_8 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 9)) begin
        _saxi_register_9 <= axislite_resetval_48;
        _saxi_flag_9 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 10)) begin
        _saxi_register_10 <= axislite_resetval_48;
        _saxi_flag_10 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 11)) begin
        _saxi_register_11 <= axislite_resetval_48;
        _saxi_flag_11 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 12)) begin
        _saxi_register_12 <= axislite_resetval_48;
        _saxi_flag_12 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 13)) begin
        _saxi_register_13 <= axislite_resetval_48;
        _saxi_flag_13 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 14)) begin
        _saxi_register_14 <= axislite_resetval_48;
        _saxi_flag_14 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 15)) begin
        _saxi_register_15 <= axislite_resetval_48;
        _saxi_flag_15 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 16)) begin
        _saxi_register_16 <= axislite_resetval_48;
        _saxi_flag_16 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 17)) begin
        _saxi_register_17 <= axislite_resetval_48;
        _saxi_flag_17 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 18)) begin
        _saxi_register_18 <= axislite_resetval_48;
        _saxi_flag_18 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 19)) begin
        _saxi_register_19 <= axislite_resetval_48;
        _saxi_flag_19 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 20)) begin
        _saxi_register_20 <= axislite_resetval_48;
        _saxi_flag_20 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 21)) begin
        _saxi_register_21 <= axislite_resetval_48;
        _saxi_flag_21 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 22)) begin
        _saxi_register_22 <= axislite_resetval_48;
        _saxi_flag_22 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 23)) begin
        _saxi_register_23 <= axislite_resetval_48;
        _saxi_flag_23 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 24)) begin
        _saxi_register_24 <= axislite_resetval_48;
        _saxi_flag_24 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 25)) begin
        _saxi_register_25 <= axislite_resetval_48;
        _saxi_flag_25 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 26)) begin
        _saxi_register_26 <= axislite_resetval_48;
        _saxi_flag_26 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 27)) begin
        _saxi_register_27 <= axislite_resetval_48;
        _saxi_flag_27 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 28)) begin
        _saxi_register_28 <= axislite_resetval_48;
        _saxi_flag_28 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 29)) begin
        _saxi_register_29 <= axislite_resetval_48;
        _saxi_flag_29 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 30)) begin
        _saxi_register_30 <= axislite_resetval_48;
        _saxi_flag_30 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 31)) begin
        _saxi_register_31 <= axislite_resetval_48;
        _saxi_flag_31 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 32)) begin
        _saxi_register_32 <= axislite_resetval_48;
        _saxi_flag_32 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 33)) begin
        _saxi_register_33 <= axislite_resetval_48;
        _saxi_flag_33 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 34)) begin
        _saxi_register_34 <= axislite_resetval_48;
        _saxi_flag_34 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 35)) begin
        _saxi_register_35 <= axislite_resetval_48;
        _saxi_flag_35 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 36)) begin
        _saxi_register_36 <= axislite_resetval_48;
        _saxi_flag_36 <= 0;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 0)) begin
        _saxi_register_0 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 1)) begin
        _saxi_register_1 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 2)) begin
        _saxi_register_2 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 3)) begin
        _saxi_register_3 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 4)) begin
        _saxi_register_4 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 5)) begin
        _saxi_register_5 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 6)) begin
        _saxi_register_6 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 7)) begin
        _saxi_register_7 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 8)) begin
        _saxi_register_8 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 9)) begin
        _saxi_register_9 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 10)) begin
        _saxi_register_10 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 11)) begin
        _saxi_register_11 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 12)) begin
        _saxi_register_12 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 13)) begin
        _saxi_register_13 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 14)) begin
        _saxi_register_14 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 15)) begin
        _saxi_register_15 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 16)) begin
        _saxi_register_16 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 17)) begin
        _saxi_register_17 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 18)) begin
        _saxi_register_18 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 19)) begin
        _saxi_register_19 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 20)) begin
        _saxi_register_20 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 21)) begin
        _saxi_register_21 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 22)) begin
        _saxi_register_22 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 23)) begin
        _saxi_register_23 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 24)) begin
        _saxi_register_24 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 25)) begin
        _saxi_register_25 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 26)) begin
        _saxi_register_26 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 27)) begin
        _saxi_register_27 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 28)) begin
        _saxi_register_28 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 29)) begin
        _saxi_register_29 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 30)) begin
        _saxi_register_30 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 31)) begin
        _saxi_register_31 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 32)) begin
        _saxi_register_32 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 33)) begin
        _saxi_register_33 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 34)) begin
        _saxi_register_34 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 35)) begin
        _saxi_register_35 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 36)) begin
        _saxi_register_36 <= saxi_wdata;
      end 
      if(_saxi_register_11[0] == 1) begin
        _saxi_register_11[0] <= 0;
        _saxi_register_9[0] <= 0;
      end 
      if(_saxi_register_11[1] == 1) begin
        _saxi_register_11[1] <= 0;
        _saxi_register_9[1] <= 0;
      end 
      if(_saxi_register_11[2] == 1) begin
        _saxi_register_11[2] <= 0;
        _saxi_register_9[2] <= 0;
      end 
      if(_saxi_register_11[3] == 1) begin
        _saxi_register_11[3] <= 0;
        _saxi_register_9[3] <= 0;
      end 
      if(_saxi_register_11[4] == 1) begin
        _saxi_register_11[4] <= 0;
        _saxi_register_9[4] <= 0;
      end 
      if(_saxi_register_11[5] == 1) begin
        _saxi_register_11[5] <= 0;
        _saxi_register_9[5] <= 0;
      end 
      if(_saxi_register_11[6] == 1) begin
        _saxi_register_11[6] <= 0;
        _saxi_register_9[6] <= 0;
      end 
      if(_saxi_register_11[7] == 1) begin
        _saxi_register_11[7] <= 0;
        _saxi_register_9[7] <= 0;
      end 
      if(_saxi_register_11[8] == 1) begin
        _saxi_register_11[8] <= 0;
        _saxi_register_9[8] <= 0;
      end 
      if(_saxi_register_11[9] == 1) begin
        _saxi_register_11[9] <= 0;
        _saxi_register_9[9] <= 0;
      end 
      if(_saxi_register_11[10] == 1) begin
        _saxi_register_11[10] <= 0;
        _saxi_register_9[10] <= 0;
      end 
      if(_saxi_register_11[11] == 1) begin
        _saxi_register_11[11] <= 0;
        _saxi_register_9[11] <= 0;
      end 
      if(_saxi_register_11[12] == 1) begin
        _saxi_register_11[12] <= 0;
        _saxi_register_9[12] <= 0;
      end 
      if(_saxi_register_11[13] == 1) begin
        _saxi_register_11[13] <= 0;
        _saxi_register_9[13] <= 0;
      end 
      if(_saxi_register_11[14] == 1) begin
        _saxi_register_11[14] <= 0;
        _saxi_register_9[14] <= 0;
      end 
      if(_saxi_register_11[15] == 1) begin
        _saxi_register_11[15] <= 0;
        _saxi_register_9[15] <= 0;
      end 
      if(_saxi_register_11[16] == 1) begin
        _saxi_register_11[16] <= 0;
        _saxi_register_9[16] <= 0;
      end 
      if(_saxi_register_11[17] == 1) begin
        _saxi_register_11[17] <= 0;
        _saxi_register_9[17] <= 0;
      end 
      if(_saxi_register_11[18] == 1) begin
        _saxi_register_11[18] <= 0;
        _saxi_register_9[18] <= 0;
      end 
      if(_saxi_register_11[19] == 1) begin
        _saxi_register_11[19] <= 0;
        _saxi_register_9[19] <= 0;
      end 
      if(_saxi_register_11[20] == 1) begin
        _saxi_register_11[20] <= 0;
        _saxi_register_9[20] <= 0;
      end 
      if(_saxi_register_11[21] == 1) begin
        _saxi_register_11[21] <= 0;
        _saxi_register_9[21] <= 0;
      end 
      if(_saxi_register_11[22] == 1) begin
        _saxi_register_11[22] <= 0;
        _saxi_register_9[22] <= 0;
      end 
      if(_saxi_register_11[23] == 1) begin
        _saxi_register_11[23] <= 0;
        _saxi_register_9[23] <= 0;
      end 
      if(_saxi_register_11[24] == 1) begin
        _saxi_register_11[24] <= 0;
        _saxi_register_9[24] <= 0;
      end 
      if(_saxi_register_11[25] == 1) begin
        _saxi_register_11[25] <= 0;
        _saxi_register_9[25] <= 0;
      end 
      if(_saxi_register_11[26] == 1) begin
        _saxi_register_11[26] <= 0;
        _saxi_register_9[26] <= 0;
      end 
      if(_saxi_register_11[27] == 1) begin
        _saxi_register_11[27] <= 0;
        _saxi_register_9[27] <= 0;
      end 
      if(_saxi_register_11[28] == 1) begin
        _saxi_register_11[28] <= 0;
        _saxi_register_9[28] <= 0;
      end 
      if(_saxi_register_11[29] == 1) begin
        _saxi_register_11[29] <= 0;
        _saxi_register_9[29] <= 0;
      end 
      if(_saxi_register_11[30] == 1) begin
        _saxi_register_11[30] <= 0;
        _saxi_register_9[30] <= 0;
      end 
      if(_saxi_register_11[31] == 1) begin
        _saxi_register_11[31] <= 0;
        _saxi_register_9[31] <= 0;
      end 
      if(irq_busy_edge_51) begin
        _saxi_register_9[0] <= irq_busy_edge_51;
      end 
      if(irq_extern_edge_53) begin
        _saxi_register_9[1] <= irq_extern_edge_53;
      end 
      if(main_fsm == 0) begin
        _saxi_register_5 <= 0;
        _saxi_register_6 <= 0;
        _saxi_register_7 <= 0;
      end 
      if(main_fsm == 1) begin
        internal_state_counter <= 0;
        _saxi_register_12 <= 0;
      end else if(main_fsm == _saxi_register_13) begin
        if(internal_state_counter == _saxi_register_14) begin
          internal_state_counter <= 0;
          _saxi_register_12 <= _saxi_register_12 + 1;
        end else begin
          internal_state_counter <= internal_state_counter + 1;
        end
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_0 <= 1;
        _saxi_flag_0 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_1 <= 1;
        _saxi_flag_1 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_2 <= 1;
        _saxi_flag_2 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_3 <= 1;
        _saxi_flag_3 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_4 <= 1;
        _saxi_flag_4 <= 0;
      end 
      if((main_fsm == 1) && 1) begin
        _saxi_register_5 <= 1;
        _saxi_flag_5 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_6 <= 1;
        _saxi_flag_6 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_7 <= 1;
        _saxi_flag_7 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_8 <= 1;
        _saxi_flag_8 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_9 <= 1;
        _saxi_flag_9 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_10 <= 1;
        _saxi_flag_10 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_11 <= 1;
        _saxi_flag_11 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_12 <= 1;
        _saxi_flag_12 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_13 <= 1;
        _saxi_flag_13 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_14 <= 1;
        _saxi_flag_14 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_15 <= 1;
        _saxi_flag_15 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_16 <= 1;
        _saxi_flag_16 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_17 <= 1;
        _saxi_flag_17 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_18 <= 1;
        _saxi_flag_18 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_19 <= 1;
        _saxi_flag_19 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_20 <= 1;
        _saxi_flag_20 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_21 <= 1;
        _saxi_flag_21 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_22 <= 1;
        _saxi_flag_22 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_23 <= 1;
        _saxi_flag_23 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_24 <= 1;
        _saxi_flag_24 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_25 <= 1;
        _saxi_flag_25 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_26 <= 1;
        _saxi_flag_26 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_27 <= 1;
        _saxi_flag_27 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_28 <= 1;
        _saxi_flag_28 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_29 <= 1;
        _saxi_flag_29 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_30 <= 1;
        _saxi_flag_30 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_31 <= 1;
        _saxi_flag_31 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_32 <= 1;
        _saxi_flag_32 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_33 <= 1;
        _saxi_flag_33 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_34 <= 1;
        _saxi_flag_34 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_35 <= 1;
        _saxi_flag_35 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_36 <= 1;
        _saxi_flag_36 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_0 <= 0;
        _saxi_flag_0 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_1 <= 0;
        _saxi_flag_1 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_2 <= 0;
        _saxi_flag_2 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_3 <= 0;
        _saxi_flag_3 <= 0;
      end 
      if((main_fsm == 2) && 1) begin
        _saxi_register_4 <= 0;
        _saxi_flag_4 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_5 <= 0;
        _saxi_flag_5 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_6 <= 0;
        _saxi_flag_6 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_7 <= 0;
        _saxi_flag_7 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_8 <= 0;
        _saxi_flag_8 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_9 <= 0;
        _saxi_flag_9 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_10 <= 0;
        _saxi_flag_10 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_11 <= 0;
        _saxi_flag_11 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_12 <= 0;
        _saxi_flag_12 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_13 <= 0;
        _saxi_flag_13 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_14 <= 0;
        _saxi_flag_14 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_15 <= 0;
        _saxi_flag_15 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_16 <= 0;
        _saxi_flag_16 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_17 <= 0;
        _saxi_flag_17 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_18 <= 0;
        _saxi_flag_18 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_19 <= 0;
        _saxi_flag_19 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_20 <= 0;
        _saxi_flag_20 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_21 <= 0;
        _saxi_flag_21 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_22 <= 0;
        _saxi_flag_22 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_23 <= 0;
        _saxi_flag_23 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_24 <= 0;
        _saxi_flag_24 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_25 <= 0;
        _saxi_flag_25 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_26 <= 0;
        _saxi_flag_26 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_27 <= 0;
        _saxi_flag_27 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_28 <= 0;
        _saxi_flag_28 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_29 <= 0;
        _saxi_flag_29 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_30 <= 0;
        _saxi_flag_30 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_31 <= 0;
        _saxi_flag_31 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_32 <= 0;
        _saxi_flag_32 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_33 <= 0;
        _saxi_flag_33 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_34 <= 0;
        _saxi_flag_34 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_35 <= 0;
        _saxi_flag_35 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_36 <= 0;
        _saxi_flag_36 <= 0;
      end 
      if((main_fsm == 159) && 0) begin
        _saxi_register_0 <= 0;
        _saxi_flag_0 <= 0;
      end 
      if((main_fsm == 159) && 0) begin
        _saxi_register_1 <= 0;
        _saxi_flag_1 <= 0;
      end 
      if((main_fsm == 159) && 0) begin
        _saxi_register_2 <= 0;
        _saxi_flag_2 <= 0;
      end 
      if((main_fsm == 159) && 0) begin
        _saxi_register_3 <= 0;
        _saxi_flag_3 <= 0;
      end 
      if((main_fsm == 159) && 0) begin
        _saxi_register_4 <= 0;
        _saxi_flag_4 <= 0;
      end 
      if((main_fsm == 159) && 1) begin
        _saxi_register_5 <= 0;
        _saxi_flag_5 <= 0;
      end 
      if((main_fsm == 159) && 0) begin
        _saxi_register_6 <= 0;
        _saxi_flag_6 <= 0;
      end 
      if((main_fsm == 159) && 0) begin
        _saxi_register_7 <= 0;
        _saxi_flag_7 <= 0;
      end 
      if((main_fsm == 159) && 0) begin
        _saxi_register_8 <= 0;
        _saxi_flag_8 <= 0;
      end 
      if((main_fsm == 159) && 0) begin
        _saxi_register_9 <= 0;
        _saxi_flag_9 <= 0;
      end 
      if((main_fsm == 159) && 0) begin
        _saxi_register_10 <= 0;
        _saxi_flag_10 <= 0;
      end 
      if((main_fsm == 159) && 0) begin
        _saxi_register_11 <= 0;
        _saxi_flag_11 <= 0;
      end 
      if((main_fsm == 159) && 0) begin
        _saxi_register_12 <= 0;
        _saxi_flag_12 <= 0;
      end 
      if((main_fsm == 159) && 0) begin
        _saxi_register_13 <= 0;
        _saxi_flag_13 <= 0;
      end 
      if((main_fsm == 159) && 0) begin
        _saxi_register_14 <= 0;
        _saxi_flag_14 <= 0;
      end 
      if((main_fsm == 159) && 0) begin
        _saxi_register_15 <= 0;
        _saxi_flag_15 <= 0;
      end 
      if((main_fsm == 159) && 0) begin
        _saxi_register_16 <= 0;
        _saxi_flag_16 <= 0;
      end 
      if((main_fsm == 159) && 0) begin
        _saxi_register_17 <= 0;
        _saxi_flag_17 <= 0;
      end 
      if((main_fsm == 159) && 0) begin
        _saxi_register_18 <= 0;
        _saxi_flag_18 <= 0;
      end 
      if((main_fsm == 159) && 0) begin
        _saxi_register_19 <= 0;
        _saxi_flag_19 <= 0;
      end 
      if((main_fsm == 159) && 0) begin
        _saxi_register_20 <= 0;
        _saxi_flag_20 <= 0;
      end 
      if((main_fsm == 159) && 0) begin
        _saxi_register_21 <= 0;
        _saxi_flag_21 <= 0;
      end 
      if((main_fsm == 159) && 0) begin
        _saxi_register_22 <= 0;
        _saxi_flag_22 <= 0;
      end 
      if((main_fsm == 159) && 0) begin
        _saxi_register_23 <= 0;
        _saxi_flag_23 <= 0;
      end 
      if((main_fsm == 159) && 0) begin
        _saxi_register_24 <= 0;
        _saxi_flag_24 <= 0;
      end 
      if((main_fsm == 159) && 0) begin
        _saxi_register_25 <= 0;
        _saxi_flag_25 <= 0;
      end 
      if((main_fsm == 159) && 0) begin
        _saxi_register_26 <= 0;
        _saxi_flag_26 <= 0;
      end 
      if((main_fsm == 159) && 0) begin
        _saxi_register_27 <= 0;
        _saxi_flag_27 <= 0;
      end 
      if((main_fsm == 159) && 0) begin
        _saxi_register_28 <= 0;
        _saxi_flag_28 <= 0;
      end 
      if((main_fsm == 159) && 0) begin
        _saxi_register_29 <= 0;
        _saxi_flag_29 <= 0;
      end 
      if((main_fsm == 159) && 0) begin
        _saxi_register_30 <= 0;
        _saxi_flag_30 <= 0;
      end 
      if((main_fsm == 159) && 0) begin
        _saxi_register_31 <= 0;
        _saxi_flag_31 <= 0;
      end 
      if((main_fsm == 159) && 0) begin
        _saxi_register_32 <= 0;
        _saxi_flag_32 <= 0;
      end 
      if((main_fsm == 159) && 0) begin
        _saxi_register_33 <= 0;
        _saxi_flag_33 <= 0;
      end 
      if((main_fsm == 159) && 0) begin
        _saxi_register_34 <= 0;
        _saxi_flag_34 <= 0;
      end 
      if((main_fsm == 159) && 0) begin
        _saxi_register_35 <= 0;
        _saxi_flag_35 <= 0;
      end 
      if((main_fsm == 159) && 0) begin
        _saxi_register_36 <= 0;
        _saxi_flag_36 <= 0;
      end 
    end
  end

  localparam _saxi_register_fsm_1 = 1;
  localparam _saxi_register_fsm_2 = 2;
  localparam _saxi_register_fsm_3 = 3;
  localparam _saxi_register_fsm_4 = 4;

  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      _saxi_register_fsm <= _saxi_register_fsm_init;
      axis_maskaddr_45 <= 0;
    end else begin
      case(_saxi_register_fsm)
        _saxi_register_fsm_init: begin
          if(readvalid_42 || writevalid_41) begin
            axis_maskaddr_45 <= (addr_40 >> _saxi_shift) & _saxi_mask;
          end 
          if(readvalid_42) begin
            _saxi_register_fsm <= _saxi_register_fsm_1;
          end 
          if(writevalid_41) begin
            _saxi_register_fsm <= _saxi_register_fsm_3;
          end 
        end
        _saxi_register_fsm_1: begin
          if(saxi_rready || !saxi_rvalid) begin
            _saxi_register_fsm <= _saxi_register_fsm_2;
          end 
        end
        _saxi_register_fsm_2: begin
          if(saxi_rready && saxi_rvalid) begin
            _saxi_register_fsm <= _saxi_register_fsm_init;
          end 
        end
        _saxi_register_fsm_3: begin
          if(saxi_wvalid) begin
            _saxi_register_fsm <= _saxi_register_fsm_4;
          end 
        end
        _saxi_register_fsm_4: begin
          if(saxi_bready && saxi_bvalid) begin
            _saxi_register_fsm <= _saxi_register_fsm_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    _rst_logic_1 <= rst_logic;
    _rst_logic_2 <= _rst_logic_1;
    RST <= rst_logic | _rst_logic_1 | _rst_logic_2;
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      irq <= 0;
    end else begin
      irq <= |irq_49;
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      irq_busy_edge_50 <= 0;
    end else begin
      irq_busy_edge_50 <= irq_busy;
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      irq_extern_edge_52 <= 0;
    end else begin
      irq_extern_edge_52 <= irq_extern;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1355_1 <= 0;
      __tmp_1706_1 <= 0;
    end else begin
      __tmp_1355_1 <= _tmp_1355;
      __tmp_1706_1 <= _tmp_1706;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1357_1 <= 0;
      __tmp_1708_1 <= 0;
    end else begin
      __tmp_1357_1 <= _tmp_1357;
      __tmp_1708_1 <= _tmp_1708;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1359_1 <= 0;
      __tmp_1710_1 <= 0;
    end else begin
      __tmp_1359_1 <= _tmp_1359;
      __tmp_1710_1 <= _tmp_1710;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1361_1 <= 0;
      __tmp_1712_1 <= 0;
    end else begin
      __tmp_1361_1 <= _tmp_1361;
      __tmp_1712_1 <= _tmp_1712;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1693_1 <= 0;
    end else begin
      __tmp_1693_1 <= _tmp_1693;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1695_1 <= 0;
    end else begin
      __tmp_1695_1 <= _tmp_1695;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1697_1 <= 0;
    end else begin
      __tmp_1697_1 <= _tmp_1697;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1699_1 <= 0;
    end else begin
      __tmp_1699_1 <= _tmp_1699;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_434_1 <= 0;
      __tmp_1460_1 <= 0;
      __tmp_1498_1 <= 0;
    end else begin
      __tmp_434_1 <= _tmp_434;
      __tmp_1460_1 <= _tmp_1460;
      __tmp_1498_1 <= _tmp_1498;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_436_1 <= 0;
      __tmp_1464_1 <= 0;
      __tmp_1500_1 <= 0;
    end else begin
      __tmp_436_1 <= _tmp_436;
      __tmp_1464_1 <= _tmp_1464;
      __tmp_1500_1 <= _tmp_1500;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_438_1 <= 0;
      __tmp_1468_1 <= 0;
      __tmp_1502_1 <= 0;
    end else begin
      __tmp_438_1 <= _tmp_438;
      __tmp_1468_1 <= _tmp_1468;
      __tmp_1502_1 <= _tmp_1502;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_440_1 <= 0;
      __tmp_1472_1 <= 0;
      __tmp_1504_1 <= 0;
    end else begin
      __tmp_440_1 <= _tmp_440;
      __tmp_1472_1 <= _tmp_1472;
      __tmp_1504_1 <= _tmp_1504;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_447_1 <= 0;
      __tmp_1612_1 <= 0;
    end else begin
      __tmp_447_1 <= _tmp_447;
      __tmp_1612_1 <= _tmp_1612;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_449_1 <= 0;
      __tmp_1616_1 <= 0;
    end else begin
      __tmp_449_1 <= _tmp_449;
      __tmp_1616_1 <= _tmp_1616;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_451_1 <= 0;
      __tmp_1620_1 <= 0;
    end else begin
      __tmp_451_1 <= _tmp_451;
      __tmp_1620_1 <= _tmp_1620;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_453_1 <= 0;
      __tmp_1624_1 <= 0;
    end else begin
      __tmp_453_1 <= _tmp_453;
      __tmp_1624_1 <= _tmp_1624;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_460_1 <= 0;
    end else begin
      __tmp_460_1 <= _tmp_460;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_462_1 <= 0;
    end else begin
      __tmp_462_1 <= _tmp_462;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_464_1 <= 0;
    end else begin
      __tmp_464_1 <= _tmp_464;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_466_1 <= 0;
    end else begin
      __tmp_466_1 <= _tmp_466;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_473_1 <= 0;
    end else begin
      __tmp_473_1 <= _tmp_473;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_475_1 <= 0;
    end else begin
      __tmp_475_1 <= _tmp_475;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_477_1 <= 0;
    end else begin
      __tmp_477_1 <= _tmp_477;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_479_1 <= 0;
    end else begin
      __tmp_479_1 <= _tmp_479;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_486_1 <= 0;
    end else begin
      __tmp_486_1 <= _tmp_486;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_488_1 <= 0;
    end else begin
      __tmp_488_1 <= _tmp_488;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_490_1 <= 0;
    end else begin
      __tmp_490_1 <= _tmp_490;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_492_1 <= 0;
    end else begin
      __tmp_492_1 <= _tmp_492;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_499_1 <= 0;
    end else begin
      __tmp_499_1 <= _tmp_499;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_501_1 <= 0;
    end else begin
      __tmp_501_1 <= _tmp_501;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_503_1 <= 0;
    end else begin
      __tmp_503_1 <= _tmp_503;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_505_1 <= 0;
    end else begin
      __tmp_505_1 <= _tmp_505;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_512_1 <= 0;
    end else begin
      __tmp_512_1 <= _tmp_512;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_514_1 <= 0;
    end else begin
      __tmp_514_1 <= _tmp_514;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_516_1 <= 0;
    end else begin
      __tmp_516_1 <= _tmp_516;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_518_1 <= 0;
    end else begin
      __tmp_518_1 <= _tmp_518;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_525_1 <= 0;
    end else begin
      __tmp_525_1 <= _tmp_525;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_527_1 <= 0;
    end else begin
      __tmp_527_1 <= _tmp_527;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_529_1 <= 0;
    end else begin
      __tmp_529_1 <= _tmp_529;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_531_1 <= 0;
    end else begin
      __tmp_531_1 <= _tmp_531;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_538_1 <= 0;
    end else begin
      __tmp_538_1 <= _tmp_538;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_540_1 <= 0;
    end else begin
      __tmp_540_1 <= _tmp_540;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_542_1 <= 0;
    end else begin
      __tmp_542_1 <= _tmp_542;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_544_1 <= 0;
    end else begin
      __tmp_544_1 <= _tmp_544;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_405_1 <= 0;
      __tmp_1664_1 <= 0;
    end else begin
      __tmp_405_1 <= _tmp_405;
      __tmp_1664_1 <= _tmp_1664;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_551_1 <= 0;
    end else begin
      __tmp_551_1 <= _tmp_551;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_553_1 <= 0;
    end else begin
      __tmp_553_1 <= _tmp_553;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_555_1 <= 0;
    end else begin
      __tmp_555_1 <= _tmp_555;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_557_1 <= 0;
    end else begin
      __tmp_557_1 <= _tmp_557;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_564_1 <= 0;
    end else begin
      __tmp_564_1 <= _tmp_564;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_566_1 <= 0;
    end else begin
      __tmp_566_1 <= _tmp_566;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_568_1 <= 0;
    end else begin
      __tmp_568_1 <= _tmp_568;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_570_1 <= 0;
    end else begin
      __tmp_570_1 <= _tmp_570;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_577_1 <= 0;
    end else begin
      __tmp_577_1 <= _tmp_577;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_579_1 <= 0;
    end else begin
      __tmp_579_1 <= _tmp_579;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_581_1 <= 0;
    end else begin
      __tmp_581_1 <= _tmp_581;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_583_1 <= 0;
    end else begin
      __tmp_583_1 <= _tmp_583;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_590_1 <= 0;
    end else begin
      __tmp_590_1 <= _tmp_590;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_592_1 <= 0;
    end else begin
      __tmp_592_1 <= _tmp_592;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_594_1 <= 0;
    end else begin
      __tmp_594_1 <= _tmp_594;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_596_1 <= 0;
    end else begin
      __tmp_596_1 <= _tmp_596;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_603_1 <= 0;
    end else begin
      __tmp_603_1 <= _tmp_603;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_605_1 <= 0;
    end else begin
      __tmp_605_1 <= _tmp_605;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_607_1 <= 0;
    end else begin
      __tmp_607_1 <= _tmp_607;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_609_1 <= 0;
    end else begin
      __tmp_609_1 <= _tmp_609;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_616_1 <= 0;
    end else begin
      __tmp_616_1 <= _tmp_616;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_618_1 <= 0;
    end else begin
      __tmp_618_1 <= _tmp_618;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_620_1 <= 0;
    end else begin
      __tmp_620_1 <= _tmp_620;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_622_1 <= 0;
    end else begin
      __tmp_622_1 <= _tmp_622;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_629_1 <= 0;
    end else begin
      __tmp_629_1 <= _tmp_629;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_631_1 <= 0;
    end else begin
      __tmp_631_1 <= _tmp_631;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_633_1 <= 0;
    end else begin
      __tmp_633_1 <= _tmp_633;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_635_1 <= 0;
    end else begin
      __tmp_635_1 <= _tmp_635;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_642_1 <= 0;
    end else begin
      __tmp_642_1 <= _tmp_642;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_644_1 <= 0;
    end else begin
      __tmp_644_1 <= _tmp_644;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_646_1 <= 0;
    end else begin
      __tmp_646_1 <= _tmp_646;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_648_1 <= 0;
    end else begin
      __tmp_648_1 <= _tmp_648;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_655_1 <= 0;
    end else begin
      __tmp_655_1 <= _tmp_655;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_657_1 <= 0;
    end else begin
      __tmp_657_1 <= _tmp_657;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_659_1 <= 0;
    end else begin
      __tmp_659_1 <= _tmp_659;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_661_1 <= 0;
    end else begin
      __tmp_661_1 <= _tmp_661;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_411_1 <= 0;
      __tmp_1670_1 <= 0;
    end else begin
      __tmp_411_1 <= _tmp_411;
      __tmp_1670_1 <= _tmp_1670;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_413_1 <= 0;
      __tmp_1672_1 <= 0;
    end else begin
      __tmp_413_1 <= _tmp_413;
      __tmp_1672_1 <= _tmp_1672;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_415_1 <= 0;
      __tmp_1674_1 <= 0;
    end else begin
      __tmp_415_1 <= _tmp_415;
      __tmp_1674_1 <= _tmp_1674;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_417_1 <= 0;
      __tmp_1676_1 <= 0;
    end else begin
      __tmp_417_1 <= _tmp_417;
      __tmp_1676_1 <= _tmp_1676;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1312_1 <= 0;
    end else begin
      __tmp_1312_1 <= _tmp_1312;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1316_1 <= 0;
    end else begin
      __tmp_1316_1 <= _tmp_1316;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1320_1 <= 0;
    end else begin
      __tmp_1320_1 <= _tmp_1320;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1324_1 <= 0;
    end else begin
      __tmp_1324_1 <= _tmp_1324;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _acc_0_x_source_ram_renable <= 0;
      _acc_0_x_source_fifo_deq <= 0;
      _acc_0_x_idle <= 1;
      _acc_0_rshift_source_ram_renable <= 0;
      _acc_0_rshift_source_fifo_deq <= 0;
      _acc_0_rshift_idle <= 1;
      _acc_0_sum_sink_wenable <= 0;
      _acc_0_sum_sink_fifo_enq <= 0;
      _acc_0_valid_sink_wenable <= 0;
      _acc_0_valid_sink_fifo_enq <= 0;
      __acc_0_stream_ivalid_1 <= 0;
      __acc_0_stream_ivalid_2 <= 0;
      _reduceadd_data_4 <= 1'sd0;
      _reduceadd_count_4 <= 0;
      _reduceadd_prev_count_max_4 <= 0;
      _pulse_data_6 <= 1'sd0;
      _pulse_count_6 <= 0;
      _pulse_prev_count_max_6 <= 0;
      __delay_data_928_sll_16 <= 0;
      __delay_data_929__variable_1 <= 0;
      __delay_data_930_eq_34 <= 0;
      _cond_data_35 <= 0;
      __delay_data_931_pulse_6 <= 0;
      __variable_wdata_3 <= 0;
      __variable_wdata_0 <= 0;
      __variable_wdata_2 <= 0;
      __variable_wdata_1 <= 0;
      _tmp_1536 <= 0;
      _tmp_1537 <= 0;
      _tmp_1538 <= 0;
      _tmp_1539 <= 0;
      _tmp_1540 <= 0;
      _tmp_1541 <= 0;
      _tmp_1542 <= 0;
      _tmp_1543 <= 0;
      _tmp_1544 <= 0;
      _tmp_1545 <= 0;
      _tmp_1546 <= 0;
      _tmp_1547 <= 0;
      _tmp_1548 <= 0;
      _tmp_1549 <= 0;
      _tmp_1550 <= 0;
      _tmp_1551 <= 0;
      _tmp_1552 <= 0;
      _tmp_1553 <= 0;
      _tmp_1554 <= 0;
      _tmp_1555 <= 0;
      _tmp_1556 <= 0;
      _tmp_1557 <= 0;
      _tmp_1558 <= 0;
      _acc_0_busy_reg <= 0;
    end else begin
      if(_acc_0_stream_oready) begin
        _acc_0_x_source_ram_renable <= 0;
        _acc_0_x_source_fifo_deq <= 0;
      end 
      _acc_0_x_idle <= _acc_0_x_idle;
      if(_acc_0_stream_oready) begin
        _acc_0_rshift_source_ram_renable <= 0;
        _acc_0_rshift_source_fifo_deq <= 0;
      end 
      _acc_0_rshift_idle <= _acc_0_rshift_idle;
      if(_acc_0_stream_oready) begin
        _acc_0_sum_sink_wenable <= 0;
        _acc_0_sum_sink_fifo_enq <= 0;
      end 
      if(_acc_0_stream_oready) begin
        _acc_0_valid_sink_wenable <= 0;
        _acc_0_valid_sink_fifo_enq <= 0;
      end 
      if(_acc_0_stream_oready) begin
        __acc_0_stream_ivalid_1 <= _acc_0_stream_ivalid;
      end 
      if(_acc_0_stream_oready) begin
        __acc_0_stream_ivalid_2 <= __acc_0_stream_ivalid_1;
      end 
      if(_acc_0_stream_ivalid && _acc_0_stream_oready && _reduceadd_reset_cond_4) begin
        _reduceadd_data_4 <= 1'sd0;
      end 
      if(_acc_0_stream_ivalid && _acc_0_stream_oready) begin
        _reduceadd_count_4 <= (_reduceadd_current_count_4 >= acc_0_size_data - 1)? 0 : _reduceadd_current_count_4 + 1;
      end 
      if(_acc_0_stream_ivalid && _acc_0_stream_oready) begin
        _reduceadd_prev_count_max_4 <= _reduceadd_current_count_4 >= acc_0_size_data - 1;
      end 
      if(_acc_0_stream_ivalid && _acc_0_stream_oready) begin
        _reduceadd_data_4 <= _reduceadd_current_data_4 + acc_0_x_data;
      end 
      if(_acc_0_stream_ivalid && _acc_0_stream_oready && _pulse_reset_cond_6) begin
        _pulse_data_6 <= 1'sd0;
      end 
      if(_acc_0_stream_ivalid && _acc_0_stream_oready) begin
        _pulse_count_6 <= (_pulse_current_count_6 >= acc_0_size_data - 1)? 0 : _pulse_current_count_6 + 1;
      end 
      if(_acc_0_stream_ivalid && _acc_0_stream_oready) begin
        _pulse_prev_count_max_6 <= _pulse_current_count_6 >= acc_0_size_data - 1;
      end 
      if(_acc_0_stream_ivalid && _acc_0_stream_oready) begin
        _pulse_data_6 <= _pulse_current_count_6 >= acc_0_size_data - 1;
      end 
      if(_acc_0_stream_oready) begin
        __delay_data_928_sll_16 <= _sll_data_16;
      end 
      if(_acc_0_stream_oready) begin
        __delay_data_929__variable_1 <= acc_0_rshift_data;
      end 
      if(_acc_0_stream_oready) begin
        __delay_data_930_eq_34 <= _eq_data_34;
      end 
      if(_acc_0_stream_oready) begin
        _cond_data_35 <= (__delay_data_930_eq_34)? _reduceadd_data_4 : _sra_data_32;
      end 
      if(_acc_0_stream_oready) begin
        __delay_data_931_pulse_6 <= _pulse_data_6;
      end 
      if(__stream_avg_pool_serial_52_stream_ivalid_3 && _stream_avg_pool_serial_52_stream_oready) begin
        __variable_wdata_3 <= __delay_data_1188__delay_1187__delay_1186__variable_915;
      end 
      if(__stream_avg_pool_serial_52_stream_ivalid_3 && _stream_avg_pool_serial_52_stream_oready) begin
        __variable_wdata_0 <= _cond_data_926;
      end 
      if(__stream_avg_pool_serial_52_stream_ivalid_3 && _stream_avg_pool_serial_52_stream_oready) begin
        __variable_wdata_2 <= __delay_data_1191__delay_1190__delay_1189__variable_912;
      end 
      if(__stream_avg_pool_serial_52_stream_ivalid_3 && _stream_avg_pool_serial_52_stream_oready) begin
        __variable_wdata_1 <= 1'sd0;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_1536 <= _acc_0_source_start;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_1537 <= _tmp_1536;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_1538 <= _tmp_1537;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_1539 <= _acc_0_source_start;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_1540 <= _tmp_1539;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_1541 <= _tmp_1540;
      end 
      if(_acc_0_stream_oready && _tmp_1541) begin
        __variable_wdata_3 <= 1;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_1542 <= _acc_0_source_start;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_1543 <= _tmp_1542;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_1544 <= _tmp_1543;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_1545 <= _tmp_1544;
      end 
      if(_acc_0_stream_oready && _tmp_1545) begin
        __variable_wdata_3 <= 0;
      end 
      if(_acc_0_stream_oready && 1'd0) begin
        __variable_wdata_3 <= 1;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_1546 <= _acc_0_source_start;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_1547 <= _tmp_1546;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_1548 <= _tmp_1547;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_1549 <= _tmp_1548;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_1550 <= _acc_0_source_stop;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_1551 <= _tmp_1550;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_1552 <= _tmp_1551;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_1553 <= _tmp_1552;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_1554 <= _acc_0_source_busy;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_1555 <= _tmp_1554;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_1556 <= _tmp_1555;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_1557 <= _tmp_1556;
      end 
      if(_acc_0_stream_oready) begin
        _tmp_1558 <= _acc_0_sink_busy;
      end 
      if(!_acc_0_sink_busy && _tmp_1558) begin
        _acc_0_busy_reg <= 0;
      end 
      if(_acc_0_source_busy) begin
        _acc_0_busy_reg <= 1;
      end 
    end
  end

  localparam _acc_0_fsm_1 = 1;
  localparam _acc_0_fsm_2 = 2;
  localparam _acc_0_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _acc_0_fsm <= _acc_0_fsm_init;
      _acc_0_source_start <= 0;
      _acc_0_source_busy <= 0;
      _acc_0_stream_ivalid <= 0;
    end else begin
      if(__stream_avg_pool_serial_52_stream_ivalid_3 && _stream_avg_pool_serial_52_stream_oready) begin
        _acc_0_stream_ivalid <= 1'd1;
      end 
      if(_stream_avg_pool_serial_52_stream_oready && _stream_avg_pool_serial_52_busy) begin
        _acc_0_source_busy <= _stream_avg_pool_serial_52_source_busy;
      end 
      if(_acc_0_stream_oready && _tmp_1538) begin
        _acc_0_stream_ivalid <= 1;
      end 
      if(_acc_0_stream_oready && 1'd0) begin
        _acc_0_stream_ivalid <= 0;
      end 
      case(_acc_0_fsm)
        _acc_0_fsm_init: begin
          if(_acc_0_run_flag) begin
            _acc_0_source_start <= 1;
          end 
          if(_acc_0_run_flag) begin
            _acc_0_fsm <= _acc_0_fsm_1;
          end 
        end
        _acc_0_fsm_1: begin
          if(_acc_0_source_start && _acc_0_stream_oready) begin
            _acc_0_source_start <= 0;
            _acc_0_source_busy <= 1;
          end 
          if(_acc_0_source_start && _acc_0_stream_oready) begin
            _acc_0_fsm <= _acc_0_fsm_2;
          end 
        end
        _acc_0_fsm_2: begin
          if(_acc_0_stream_oready) begin
            _acc_0_fsm <= _acc_0_fsm_3;
          end 
        end
        _acc_0_fsm_3: begin
          if(_acc_0_stream_oready && 1'd0) begin
            _acc_0_source_busy <= 0;
          end 
          if(_acc_0_stream_oready && 1'd0 && _acc_0_run_flag) begin
            _acc_0_source_start <= 1;
          end 
          if(_acc_0_stream_oready && 1'd0) begin
            _acc_0_fsm <= _acc_0_fsm_init;
          end 
          if(_acc_0_stream_oready && 1'd0 && _acc_0_run_flag) begin
            _acc_0_fsm <= _acc_0_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _acc_1_x_source_ram_renable <= 0;
      _acc_1_x_source_fifo_deq <= 0;
      _acc_1_x_idle <= 1;
      _acc_1_rshift_source_ram_renable <= 0;
      _acc_1_rshift_source_fifo_deq <= 0;
      _acc_1_rshift_idle <= 1;
      _acc_1_sum_sink_wenable <= 0;
      _acc_1_sum_sink_fifo_enq <= 0;
      _acc_1_valid_sink_wenable <= 0;
      _acc_1_valid_sink_fifo_enq <= 0;
      __acc_1_stream_ivalid_1 <= 0;
      __acc_1_stream_ivalid_2 <= 0;
      __acc_1_stream_ivalid_3 <= 0;
      __acc_1_stream_ivalid_4 <= 0;
      __acc_1_stream_ivalid_5 <= 0;
      _greaterthan_data_39 <= 0;
      _minus_data_41 <= 0;
      _reduceadd_data_52 <= 1'sd0;
      _reduceadd_count_52 <= 0;
      _reduceadd_prev_count_max_52 <= 0;
      _pulse_data_54 <= 1'sd0;
      _pulse_count_54 <= 0;
      _pulse_prev_count_max_54 <= 0;
      __delay_data_859__variable_37 <= 0;
      _sll_data_43 <= 0;
      __delay_data_856_greaterthan_39 <= 0;
      __delay_data_857_reduceadd_52 <= 0;
      __delay_data_860__delay_859__variable_37 <= 0;
      __delay_data_863_pulse_54 <= 0;
      _cond_data_49 <= 0;
      __delay_data_858__delay_857_reduceadd_52 <= 0;
      __delay_data_861__delay_860__delay_859__variable_37 <= 0;
      __delay_data_864__delay_863_pulse_54 <= 0;
      _plus_data_56 <= 0;
      __delay_data_862__delay_861__delay_860__delay_859__variable_37 <= 0;
      __delay_data_865__delay_864__delay_863_pulse_54 <= 0;
      _sra_data_57 <= 0;
      __delay_data_866__delay_865__delay_864__delay_863_pulse_54 <= 0;
      __variable_wdata_51 <= 0;
      __variable_wdata_36 <= 0;
      __variable_wdata_37 <= 0;
      __variable_wdata_38 <= 0;
      _tmp_1090 <= 0;
      _tmp_1091 <= 0;
      _tmp_1092 <= 0;
      _tmp_1093 <= 0;
      _tmp_1094 <= 0;
      _tmp_1095 <= 0;
      _tmp_1096 <= 0;
      _tmp_1097 <= 0;
      _tmp_1098 <= 0;
      _tmp_1099 <= 0;
      _tmp_1100 <= 0;
      _tmp_1101 <= 0;
      _tmp_1102 <= 0;
      _tmp_1103 <= 0;
      _tmp_1104 <= 0;
      _tmp_1105 <= 0;
      _tmp_1106 <= 0;
      _tmp_1107 <= 0;
      _tmp_1108 <= 0;
      _tmp_1109 <= 0;
      _tmp_1110 <= 0;
      _tmp_1111 <= 0;
      _tmp_1112 <= 0;
      _tmp_1113 <= 0;
      _tmp_1114 <= 0;
      _tmp_1115 <= 0;
      _tmp_1116 <= 0;
      _tmp_1117 <= 0;
      _tmp_1118 <= 0;
      _tmp_1119 <= 0;
      _tmp_1120 <= 0;
      _tmp_1121 <= 0;
      _acc_1_busy_reg <= 0;
    end else begin
      if(_acc_1_stream_oready) begin
        _acc_1_x_source_ram_renable <= 0;
        _acc_1_x_source_fifo_deq <= 0;
      end 
      _acc_1_x_idle <= _acc_1_x_idle;
      if(_acc_1_stream_oready) begin
        _acc_1_rshift_source_ram_renable <= 0;
        _acc_1_rshift_source_fifo_deq <= 0;
      end 
      _acc_1_rshift_idle <= _acc_1_rshift_idle;
      if(_acc_1_stream_oready) begin
        _acc_1_sum_sink_wenable <= 0;
        _acc_1_sum_sink_fifo_enq <= 0;
      end 
      if(_acc_1_stream_oready) begin
        _acc_1_valid_sink_wenable <= 0;
        _acc_1_valid_sink_fifo_enq <= 0;
      end 
      if(_acc_1_stream_oready) begin
        __acc_1_stream_ivalid_1 <= _acc_1_stream_ivalid;
      end 
      if(_acc_1_stream_oready) begin
        __acc_1_stream_ivalid_2 <= __acc_1_stream_ivalid_1;
      end 
      if(_acc_1_stream_oready) begin
        __acc_1_stream_ivalid_3 <= __acc_1_stream_ivalid_2;
      end 
      if(_acc_1_stream_oready) begin
        __acc_1_stream_ivalid_4 <= __acc_1_stream_ivalid_3;
      end 
      if(_acc_1_stream_oready) begin
        __acc_1_stream_ivalid_5 <= __acc_1_stream_ivalid_4;
      end 
      if(_acc_1_stream_oready) begin
        _greaterthan_data_39 <= acc_1_rshift_data > 1'sd0;
      end 
      if(_acc_1_stream_oready) begin
        _minus_data_41 <= acc_1_rshift_data - 2'sd1;
      end 
      if(_acc_1_stream_ivalid && _acc_1_stream_oready && _reduceadd_reset_cond_52) begin
        _reduceadd_data_52 <= 1'sd0;
      end 
      if(_acc_1_stream_ivalid && _acc_1_stream_oready) begin
        _reduceadd_count_52 <= (_reduceadd_current_count_52 >= acc_1_size_data - 1)? 0 : _reduceadd_current_count_52 + 1;
      end 
      if(_acc_1_stream_ivalid && _acc_1_stream_oready) begin
        _reduceadd_prev_count_max_52 <= _reduceadd_current_count_52 >= acc_1_size_data - 1;
      end 
      if(_acc_1_stream_ivalid && _acc_1_stream_oready) begin
        _reduceadd_data_52 <= _reduceadd_current_data_52 + acc_1_x_data;
      end 
      if(_acc_1_stream_ivalid && _acc_1_stream_oready && _pulse_reset_cond_54) begin
        _pulse_data_54 <= 1'sd0;
      end 
      if(_acc_1_stream_ivalid && _acc_1_stream_oready) begin
        _pulse_count_54 <= (_pulse_current_count_54 >= acc_1_size_data - 1)? 0 : _pulse_current_count_54 + 1;
      end 
      if(_acc_1_stream_ivalid && _acc_1_stream_oready) begin
        _pulse_prev_count_max_54 <= _pulse_current_count_54 >= acc_1_size_data - 1;
      end 
      if(_acc_1_stream_ivalid && _acc_1_stream_oready) begin
        _pulse_data_54 <= _pulse_current_count_54 >= acc_1_size_data - 1;
      end 
      if(_acc_1_stream_oready) begin
        __delay_data_859__variable_37 <= acc_1_rshift_data;
      end 
      if(_acc_1_stream_oready) begin
        _sll_data_43 <= 2'sd1 << _minus_data_41;
      end 
      if(_acc_1_stream_oready) begin
        __delay_data_856_greaterthan_39 <= _greaterthan_data_39;
      end 
      if(_acc_1_stream_oready) begin
        __delay_data_857_reduceadd_52 <= _reduceadd_data_52;
      end 
      if(_acc_1_stream_oready) begin
        __delay_data_860__delay_859__variable_37 <= __delay_data_859__variable_37;
      end 
      if(_acc_1_stream_oready) begin
        __delay_data_863_pulse_54 <= _pulse_data_54;
      end 
      if(_acc_1_stream_oready) begin
        _cond_data_49 <= (__delay_data_856_greaterthan_39)? _sll_data_43 : 1'sd0;
      end 
      if(_acc_1_stream_oready) begin
        __delay_data_858__delay_857_reduceadd_52 <= __delay_data_857_reduceadd_52;
      end 
      if(_acc_1_stream_oready) begin
        __delay_data_861__delay_860__delay_859__variable_37 <= __delay_data_860__delay_859__variable_37;
      end 
      if(_acc_1_stream_oready) begin
        __delay_data_864__delay_863_pulse_54 <= __delay_data_863_pulse_54;
      end 
      if(_acc_1_stream_oready) begin
        _plus_data_56 <= __delay_data_858__delay_857_reduceadd_52 + _cond_data_49;
      end 
      if(_acc_1_stream_oready) begin
        __delay_data_862__delay_861__delay_860__delay_859__variable_37 <= __delay_data_861__delay_860__delay_859__variable_37;
      end 
      if(_acc_1_stream_oready) begin
        __delay_data_865__delay_864__delay_863_pulse_54 <= __delay_data_864__delay_863_pulse_54;
      end 
      if(_acc_1_stream_oready) begin
        _sra_data_57 <= _plus_data_56 >>> __delay_data_862__delay_861__delay_860__delay_859__variable_37;
      end 
      if(_acc_1_stream_oready) begin
        __delay_data_866__delay_865__delay_864__delay_863_pulse_54 <= __delay_data_865__delay_864__delay_863_pulse_54;
      end 
      if(__stream_conv2d_24_stream_ivalid_13 && _stream_conv2d_24_stream_oready) begin
        __variable_wdata_51 <= __delay_data_1077__delay_1076__delay_1075____variable_309;
      end 
      if(__stream_conv2d_24_stream_ivalid_13 && _stream_conv2d_24_stream_oready) begin
        __variable_wdata_36 <= __substreamoutput_data_854;
      end 
      if(__stream_conv2d_24_stream_ivalid_13 && _stream_conv2d_24_stream_oready) begin
        __variable_wdata_37 <= __delay_data_1089__delay_1088__delay_1087__delay_1086___plus_867;
      end 
      if(__stream_conv2d_24_stream_ivalid_13 && _stream_conv2d_24_stream_oready) begin
        __variable_wdata_38 <= __delay_data_1102__delay_1101__delay_1100____variable_304;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1090 <= _acc_1_source_start;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1091 <= _tmp_1090;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1092 <= _tmp_1091;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1093 <= _acc_1_source_start;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1094 <= _tmp_1093;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1095 <= _tmp_1094;
      end 
      if(_acc_1_stream_oready && _tmp_1095) begin
        __variable_wdata_51 <= 1;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1096 <= _acc_1_source_start;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1097 <= _tmp_1096;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1098 <= _tmp_1097;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1099 <= _tmp_1098;
      end 
      if(_acc_1_stream_oready && _tmp_1099) begin
        __variable_wdata_51 <= 0;
      end 
      if(_acc_1_stream_oready && 1'd0) begin
        __variable_wdata_51 <= 1;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1100 <= _acc_1_source_start;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1101 <= _tmp_1100;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1102 <= _tmp_1101;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1103 <= _tmp_1102;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1104 <= _tmp_1103;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1105 <= _tmp_1104;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1106 <= _tmp_1105;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1107 <= _acc_1_source_stop;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1108 <= _tmp_1107;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1109 <= _tmp_1108;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1110 <= _tmp_1109;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1111 <= _tmp_1110;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1112 <= _tmp_1111;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1113 <= _tmp_1112;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1114 <= _acc_1_source_busy;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1115 <= _tmp_1114;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1116 <= _tmp_1115;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1117 <= _tmp_1116;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1118 <= _tmp_1117;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1119 <= _tmp_1118;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1120 <= _tmp_1119;
      end 
      if(_acc_1_stream_oready) begin
        _tmp_1121 <= _acc_1_sink_busy;
      end 
      if(!_acc_1_sink_busy && _tmp_1121) begin
        _acc_1_busy_reg <= 0;
      end 
      if(_acc_1_source_busy) begin
        _acc_1_busy_reg <= 1;
      end 
      if(__stream_matmul_55_stream_ivalid_11 && _stream_matmul_55_stream_oready) begin
        __variable_wdata_51 <= __delay_data_1205__delay_1204__delay_1203____variable_941;
      end 
      if(__stream_matmul_55_stream_ivalid_11 && _stream_matmul_55_stream_oready) begin
        __variable_wdata_36 <= __substreamoutput_data_1018;
      end 
      if(__stream_matmul_55_stream_ivalid_11 && _stream_matmul_55_stream_oready) begin
        __variable_wdata_37 <= __delay_data_1215__delay_1214__delay_1213___plus_1020;
      end 
      if(__stream_matmul_55_stream_ivalid_11 && _stream_matmul_55_stream_oready) begin
        __variable_wdata_38 <= __delay_data_1226__delay_1225__delay_1224____variable_936;
      end 
    end
  end

  localparam _acc_1_fsm_1 = 1;
  localparam _acc_1_fsm_2 = 2;
  localparam _acc_1_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _acc_1_fsm <= _acc_1_fsm_init;
      _acc_1_source_start <= 0;
      _acc_1_source_busy <= 0;
      _acc_1_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_24_stream_ivalid_13 && _stream_conv2d_24_stream_oready) begin
        _acc_1_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_24_stream_oready && _stream_conv2d_24_busy) begin
        _acc_1_source_busy <= _stream_conv2d_24_source_busy;
      end 
      if(_acc_1_stream_oready && _tmp_1092) begin
        _acc_1_stream_ivalid <= 1;
      end 
      if(_acc_1_stream_oready && 1'd0) begin
        _acc_1_stream_ivalid <= 0;
      end 
      if(__stream_matmul_55_stream_ivalid_11 && _stream_matmul_55_stream_oready) begin
        _acc_1_stream_ivalid <= 1'd1;
      end 
      if(_stream_matmul_55_stream_oready && _stream_matmul_55_busy) begin
        _acc_1_source_busy <= _stream_matmul_55_source_busy;
      end 
      case(_acc_1_fsm)
        _acc_1_fsm_init: begin
          if(_acc_1_run_flag) begin
            _acc_1_source_start <= 1;
          end 
          if(_acc_1_run_flag) begin
            _acc_1_fsm <= _acc_1_fsm_1;
          end 
        end
        _acc_1_fsm_1: begin
          if(_acc_1_source_start && _acc_1_stream_oready) begin
            _acc_1_source_start <= 0;
            _acc_1_source_busy <= 1;
          end 
          if(_acc_1_source_start && _acc_1_stream_oready) begin
            _acc_1_fsm <= _acc_1_fsm_2;
          end 
        end
        _acc_1_fsm_2: begin
          if(_acc_1_stream_oready) begin
            _acc_1_fsm <= _acc_1_fsm_3;
          end 
        end
        _acc_1_fsm_3: begin
          if(_acc_1_stream_oready && 1'd0) begin
            _acc_1_source_busy <= 0;
          end 
          if(_acc_1_stream_oready && 1'd0 && _acc_1_run_flag) begin
            _acc_1_source_start <= 1;
          end 
          if(_acc_1_stream_oready && 1'd0) begin
            _acc_1_fsm <= _acc_1_fsm_init;
          end 
          if(_acc_1_stream_oready && 1'd0 && _acc_1_run_flag) begin
            _acc_1_fsm <= _acc_1_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _add_tree_2_var0_source_ram_renable <= 0;
      _add_tree_2_var0_source_fifo_deq <= 0;
      _add_tree_2_var0_idle <= 1;
      _add_tree_2_sum_sink_wenable <= 0;
      _add_tree_2_sum_sink_fifo_enq <= 0;
      __variable_wdata_58 <= 0;
      _tmp_1813 <= 0;
      _tmp_1814 <= 0;
      _tmp_1815 <= 0;
      _tmp_1816 <= 0;
      _tmp_1817 <= 0;
      _tmp_1818 <= 0;
      _tmp_1819 <= 0;
      _tmp_1820 <= 0;
      _tmp_1821 <= 0;
      _tmp_1822 <= 0;
      _add_tree_2_busy_reg <= 0;
    end else begin
      if(_add_tree_2_stream_oready) begin
        _add_tree_2_var0_source_ram_renable <= 0;
        _add_tree_2_var0_source_fifo_deq <= 0;
      end 
      _add_tree_2_var0_idle <= _add_tree_2_var0_idle;
      if(_add_tree_2_stream_oready) begin
        _add_tree_2_sum_sink_wenable <= 0;
        _add_tree_2_sum_sink_fifo_enq <= 0;
      end 
      if(__stream_matmul_55_stream_ivalid_10 && _stream_matmul_55_stream_oready) begin
        __variable_wdata_58 <= __substreamoutput_data_1016;
      end 
      if(_add_tree_2_stream_oready) begin
        _tmp_1813 <= _add_tree_2_source_start;
      end 
      if(_add_tree_2_stream_oready) begin
        _tmp_1814 <= _tmp_1813;
      end 
      if(_add_tree_2_stream_oready) begin
        _tmp_1815 <= _tmp_1814;
      end 
      if(_add_tree_2_stream_oready) begin
        _tmp_1816 <= _add_tree_2_source_start;
      end 
      if(_add_tree_2_stream_oready) begin
        _tmp_1817 <= _tmp_1816;
      end 
      if(_add_tree_2_stream_oready) begin
        _tmp_1818 <= _add_tree_2_source_stop;
      end 
      if(_add_tree_2_stream_oready) begin
        _tmp_1819 <= _tmp_1818;
      end 
      if(_add_tree_2_stream_oready) begin
        _tmp_1820 <= _add_tree_2_source_busy;
      end 
      if(_add_tree_2_stream_oready) begin
        _tmp_1821 <= _tmp_1820;
      end 
      if(_add_tree_2_stream_oready) begin
        _tmp_1822 <= _add_tree_2_sink_busy;
      end 
      if(!_add_tree_2_sink_busy && _tmp_1822) begin
        _add_tree_2_busy_reg <= 0;
      end 
      if(_add_tree_2_source_busy) begin
        _add_tree_2_busy_reg <= 1;
      end 
    end
  end

  localparam _add_tree_2_fsm_1 = 1;
  localparam _add_tree_2_fsm_2 = 2;
  localparam _add_tree_2_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _add_tree_2_fsm <= _add_tree_2_fsm_init;
      _add_tree_2_source_start <= 0;
      _add_tree_2_source_busy <= 0;
      _add_tree_2_stream_ivalid <= 0;
    end else begin
      if(__stream_matmul_55_stream_ivalid_10 && _stream_matmul_55_stream_oready) begin
        _add_tree_2_stream_ivalid <= 1'd1;
      end 
      if(_stream_matmul_55_stream_oready && _stream_matmul_55_busy) begin
        _add_tree_2_source_busy <= _stream_matmul_55_source_busy;
      end 
      if(_add_tree_2_stream_oready && _tmp_1815) begin
        _add_tree_2_stream_ivalid <= 1;
      end 
      if(_add_tree_2_stream_oready && 1'd0) begin
        _add_tree_2_stream_ivalid <= 0;
      end 
      case(_add_tree_2_fsm)
        _add_tree_2_fsm_init: begin
          if(_add_tree_2_run_flag) begin
            _add_tree_2_source_start <= 1;
          end 
          if(_add_tree_2_run_flag) begin
            _add_tree_2_fsm <= _add_tree_2_fsm_1;
          end 
        end
        _add_tree_2_fsm_1: begin
          if(_add_tree_2_source_start && _add_tree_2_stream_oready) begin
            _add_tree_2_source_start <= 0;
            _add_tree_2_source_busy <= 1;
          end 
          if(_add_tree_2_source_start && _add_tree_2_stream_oready) begin
            _add_tree_2_fsm <= _add_tree_2_fsm_2;
          end 
        end
        _add_tree_2_fsm_2: begin
          if(_add_tree_2_stream_oready) begin
            _add_tree_2_fsm <= _add_tree_2_fsm_3;
          end 
        end
        _add_tree_2_fsm_3: begin
          if(_add_tree_2_stream_oready && 1'd0) begin
            _add_tree_2_source_busy <= 0;
          end 
          if(_add_tree_2_stream_oready && 1'd0 && _add_tree_2_run_flag) begin
            _add_tree_2_source_start <= 1;
          end 
          if(_add_tree_2_stream_oready && 1'd0) begin
            _add_tree_2_fsm <= _add_tree_2_fsm_init;
          end 
          if(_add_tree_2_stream_oready && 1'd0 && _add_tree_2_run_flag) begin
            _add_tree_2_fsm <= _add_tree_2_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _add_tree_3_var0_source_ram_renable <= 0;
      _add_tree_3_var0_source_fifo_deq <= 0;
      _add_tree_3_var0_idle <= 1;
      _add_tree_3_var1_source_ram_renable <= 0;
      _add_tree_3_var1_source_fifo_deq <= 0;
      _add_tree_3_var1_idle <= 1;
      _add_tree_3_var2_source_ram_renable <= 0;
      _add_tree_3_var2_source_fifo_deq <= 0;
      _add_tree_3_var2_idle <= 1;
      _add_tree_3_var3_source_ram_renable <= 0;
      _add_tree_3_var3_source_fifo_deq <= 0;
      _add_tree_3_var3_idle <= 1;
      _add_tree_3_var4_source_ram_renable <= 0;
      _add_tree_3_var4_source_fifo_deq <= 0;
      _add_tree_3_var4_idle <= 1;
      _add_tree_3_var5_source_ram_renable <= 0;
      _add_tree_3_var5_source_fifo_deq <= 0;
      _add_tree_3_var5_idle <= 1;
      _add_tree_3_var6_source_ram_renable <= 0;
      _add_tree_3_var6_source_fifo_deq <= 0;
      _add_tree_3_var6_idle <= 1;
      _add_tree_3_var7_source_ram_renable <= 0;
      _add_tree_3_var7_source_fifo_deq <= 0;
      _add_tree_3_var7_idle <= 1;
      _add_tree_3_var8_source_ram_renable <= 0;
      _add_tree_3_var8_source_fifo_deq <= 0;
      _add_tree_3_var8_idle <= 1;
      _add_tree_3_sum_sink_wenable <= 0;
      _add_tree_3_sum_sink_fifo_enq <= 0;
      __add_tree_3_stream_ivalid_1 <= 0;
      __add_tree_3_stream_ivalid_2 <= 0;
      __plusn_data_70 <= 0;
      __plusn_data_71 <= 0;
      __plusn_data_72 <= 0;
      __plusn_data_73 <= 0;
      __variable_wdata_60 <= 0;
      __variable_wdata_61 <= 0;
      __variable_wdata_62 <= 0;
      __variable_wdata_63 <= 0;
      __variable_wdata_64 <= 0;
      __variable_wdata_65 <= 0;
      __variable_wdata_66 <= 0;
      __variable_wdata_67 <= 0;
      __variable_wdata_68 <= 0;
      _tmp_1074 <= 0;
      _tmp_1075 <= 0;
      _tmp_1076 <= 0;
      _tmp_1077 <= 0;
      _tmp_1078 <= 0;
      _tmp_1079 <= 0;
      _tmp_1080 <= 0;
      _tmp_1081 <= 0;
      _tmp_1082 <= 0;
      _tmp_1083 <= 0;
      _tmp_1084 <= 0;
      _tmp_1085 <= 0;
      _tmp_1086 <= 0;
      _tmp_1087 <= 0;
      _tmp_1088 <= 0;
      _tmp_1089 <= 0;
      _add_tree_3_busy_reg <= 0;
    end else begin
      if(_add_tree_3_stream_oready) begin
        _add_tree_3_var0_source_ram_renable <= 0;
        _add_tree_3_var0_source_fifo_deq <= 0;
      end 
      _add_tree_3_var0_idle <= _add_tree_3_var0_idle;
      if(_add_tree_3_stream_oready) begin
        _add_tree_3_var1_source_ram_renable <= 0;
        _add_tree_3_var1_source_fifo_deq <= 0;
      end 
      _add_tree_3_var1_idle <= _add_tree_3_var1_idle;
      if(_add_tree_3_stream_oready) begin
        _add_tree_3_var2_source_ram_renable <= 0;
        _add_tree_3_var2_source_fifo_deq <= 0;
      end 
      _add_tree_3_var2_idle <= _add_tree_3_var2_idle;
      if(_add_tree_3_stream_oready) begin
        _add_tree_3_var3_source_ram_renable <= 0;
        _add_tree_3_var3_source_fifo_deq <= 0;
      end 
      _add_tree_3_var3_idle <= _add_tree_3_var3_idle;
      if(_add_tree_3_stream_oready) begin
        _add_tree_3_var4_source_ram_renable <= 0;
        _add_tree_3_var4_source_fifo_deq <= 0;
      end 
      _add_tree_3_var4_idle <= _add_tree_3_var4_idle;
      if(_add_tree_3_stream_oready) begin
        _add_tree_3_var5_source_ram_renable <= 0;
        _add_tree_3_var5_source_fifo_deq <= 0;
      end 
      _add_tree_3_var5_idle <= _add_tree_3_var5_idle;
      if(_add_tree_3_stream_oready) begin
        _add_tree_3_var6_source_ram_renable <= 0;
        _add_tree_3_var6_source_fifo_deq <= 0;
      end 
      _add_tree_3_var6_idle <= _add_tree_3_var6_idle;
      if(_add_tree_3_stream_oready) begin
        _add_tree_3_var7_source_ram_renable <= 0;
        _add_tree_3_var7_source_fifo_deq <= 0;
      end 
      _add_tree_3_var7_idle <= _add_tree_3_var7_idle;
      if(_add_tree_3_stream_oready) begin
        _add_tree_3_var8_source_ram_renable <= 0;
        _add_tree_3_var8_source_fifo_deq <= 0;
      end 
      _add_tree_3_var8_idle <= _add_tree_3_var8_idle;
      if(_add_tree_3_stream_oready) begin
        _add_tree_3_sum_sink_wenable <= 0;
        _add_tree_3_sum_sink_fifo_enq <= 0;
      end 
      if(_add_tree_3_stream_oready) begin
        __add_tree_3_stream_ivalid_1 <= _add_tree_3_stream_ivalid;
      end 
      if(_add_tree_3_stream_oready) begin
        __add_tree_3_stream_ivalid_2 <= __add_tree_3_stream_ivalid_1;
      end 
      if(_add_tree_3_stream_oready) begin
        __plusn_data_70 <= add_tree_3_var0_data + add_tree_3_var1_data + add_tree_3_var2_data;
      end 
      if(_add_tree_3_stream_oready) begin
        __plusn_data_71 <= add_tree_3_var3_data + add_tree_3_var4_data + add_tree_3_var5_data;
      end 
      if(_add_tree_3_stream_oready) begin
        __plusn_data_72 <= add_tree_3_var6_data + add_tree_3_var7_data + add_tree_3_var8_data;
      end 
      if(_add_tree_3_stream_oready) begin
        __plusn_data_73 <= __plusn_data_70 + __plusn_data_71 + __plusn_data_72;
      end 
      if(__stream_conv2d_24_stream_ivalid_10 && _stream_conv2d_24_stream_oready) begin
        __variable_wdata_60 <= __substreamoutput_data_700;
      end 
      if(__stream_conv2d_24_stream_ivalid_10 && _stream_conv2d_24_stream_oready) begin
        __variable_wdata_61 <= __substreamoutput_data_719;
      end 
      if(__stream_conv2d_24_stream_ivalid_10 && _stream_conv2d_24_stream_oready) begin
        __variable_wdata_62 <= __substreamoutput_data_738;
      end 
      if(__stream_conv2d_24_stream_ivalid_10 && _stream_conv2d_24_stream_oready) begin
        __variable_wdata_63 <= __substreamoutput_data_757;
      end 
      if(__stream_conv2d_24_stream_ivalid_10 && _stream_conv2d_24_stream_oready) begin
        __variable_wdata_64 <= __substreamoutput_data_776;
      end 
      if(__stream_conv2d_24_stream_ivalid_10 && _stream_conv2d_24_stream_oready) begin
        __variable_wdata_65 <= __substreamoutput_data_795;
      end 
      if(__stream_conv2d_24_stream_ivalid_10 && _stream_conv2d_24_stream_oready) begin
        __variable_wdata_66 <= __substreamoutput_data_814;
      end 
      if(__stream_conv2d_24_stream_ivalid_10 && _stream_conv2d_24_stream_oready) begin
        __variable_wdata_67 <= __substreamoutput_data_833;
      end 
      if(__stream_conv2d_24_stream_ivalid_10 && _stream_conv2d_24_stream_oready) begin
        __variable_wdata_68 <= __substreamoutput_data_852;
      end 
      if(_add_tree_3_stream_oready) begin
        _tmp_1074 <= _add_tree_3_source_start;
      end 
      if(_add_tree_3_stream_oready) begin
        _tmp_1075 <= _tmp_1074;
      end 
      if(_add_tree_3_stream_oready) begin
        _tmp_1076 <= _tmp_1075;
      end 
      if(_add_tree_3_stream_oready) begin
        _tmp_1077 <= _add_tree_3_source_start;
      end 
      if(_add_tree_3_stream_oready) begin
        _tmp_1078 <= _tmp_1077;
      end 
      if(_add_tree_3_stream_oready) begin
        _tmp_1079 <= _tmp_1078;
      end 
      if(_add_tree_3_stream_oready) begin
        _tmp_1080 <= _tmp_1079;
      end 
      if(_add_tree_3_stream_oready) begin
        _tmp_1081 <= _add_tree_3_source_stop;
      end 
      if(_add_tree_3_stream_oready) begin
        _tmp_1082 <= _tmp_1081;
      end 
      if(_add_tree_3_stream_oready) begin
        _tmp_1083 <= _tmp_1082;
      end 
      if(_add_tree_3_stream_oready) begin
        _tmp_1084 <= _tmp_1083;
      end 
      if(_add_tree_3_stream_oready) begin
        _tmp_1085 <= _add_tree_3_source_busy;
      end 
      if(_add_tree_3_stream_oready) begin
        _tmp_1086 <= _tmp_1085;
      end 
      if(_add_tree_3_stream_oready) begin
        _tmp_1087 <= _tmp_1086;
      end 
      if(_add_tree_3_stream_oready) begin
        _tmp_1088 <= _tmp_1087;
      end 
      if(_add_tree_3_stream_oready) begin
        _tmp_1089 <= _add_tree_3_sink_busy;
      end 
      if(!_add_tree_3_sink_busy && _tmp_1089) begin
        _add_tree_3_busy_reg <= 0;
      end 
      if(_add_tree_3_source_busy) begin
        _add_tree_3_busy_reg <= 1;
      end 
    end
  end

  localparam _add_tree_3_fsm_1 = 1;
  localparam _add_tree_3_fsm_2 = 2;
  localparam _add_tree_3_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _add_tree_3_fsm <= _add_tree_3_fsm_init;
      _add_tree_3_source_start <= 0;
      _add_tree_3_source_busy <= 0;
      _add_tree_3_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_24_stream_ivalid_10 && _stream_conv2d_24_stream_oready) begin
        _add_tree_3_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_24_stream_oready && _stream_conv2d_24_busy) begin
        _add_tree_3_source_busy <= _stream_conv2d_24_source_busy;
      end 
      if(_add_tree_3_stream_oready && _tmp_1076) begin
        _add_tree_3_stream_ivalid <= 1;
      end 
      if(_add_tree_3_stream_oready && 1'd0) begin
        _add_tree_3_stream_ivalid <= 0;
      end 
      case(_add_tree_3_fsm)
        _add_tree_3_fsm_init: begin
          if(_add_tree_3_run_flag) begin
            _add_tree_3_source_start <= 1;
          end 
          if(_add_tree_3_run_flag) begin
            _add_tree_3_fsm <= _add_tree_3_fsm_1;
          end 
        end
        _add_tree_3_fsm_1: begin
          if(_add_tree_3_source_start && _add_tree_3_stream_oready) begin
            _add_tree_3_source_start <= 0;
            _add_tree_3_source_busy <= 1;
          end 
          if(_add_tree_3_source_start && _add_tree_3_stream_oready) begin
            _add_tree_3_fsm <= _add_tree_3_fsm_2;
          end 
        end
        _add_tree_3_fsm_2: begin
          if(_add_tree_3_stream_oready) begin
            _add_tree_3_fsm <= _add_tree_3_fsm_3;
          end 
        end
        _add_tree_3_fsm_3: begin
          if(_add_tree_3_stream_oready && 1'd0) begin
            _add_tree_3_source_busy <= 0;
          end 
          if(_add_tree_3_stream_oready && 1'd0 && _add_tree_3_run_flag) begin
            _add_tree_3_source_start <= 1;
          end 
          if(_add_tree_3_stream_oready && 1'd0) begin
            _add_tree_3_fsm <= _add_tree_3_fsm_init;
          end 
          if(_add_tree_3_stream_oready && 1'd0 && _add_tree_3_run_flag) begin
            _add_tree_3_fsm <= _add_tree_3_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_rshift_round_clip_4_x_source_ram_renable <= 0;
      _mul_rshift_round_clip_4_x_source_fifo_deq <= 0;
      _mul_rshift_round_clip_4_x_idle <= 1;
      _mul_rshift_round_clip_4_y_source_ram_renable <= 0;
      _mul_rshift_round_clip_4_y_source_fifo_deq <= 0;
      _mul_rshift_round_clip_4_y_idle <= 1;
      _mul_rshift_round_clip_4_rshift_source_ram_renable <= 0;
      _mul_rshift_round_clip_4_rshift_source_fifo_deq <= 0;
      _mul_rshift_round_clip_4_rshift_idle <= 1;
      _mul_rshift_round_clip_4_z_sink_wenable <= 0;
      _mul_rshift_round_clip_4_z_sink_fifo_enq <= 0;
      __mul_rshift_round_clip_4_stream_ivalid_1 <= 0;
      __mul_rshift_round_clip_4_stream_ivalid_2 <= 0;
      __mul_rshift_round_clip_4_stream_ivalid_3 <= 0;
      __mul_rshift_round_clip_4_stream_ivalid_4 <= 0;
      __mul_rshift_round_clip_4_stream_ivalid_5 <= 0;
      __mul_rshift_round_clip_4_stream_ivalid_6 <= 0;
      __mul_rshift_round_clip_4_stream_ivalid_7 <= 0;
      __mul_rshift_round_clip_4_stream_ivalid_8 <= 0;
      _times_mul_odata_reg_77 <= 0;
      __delay_data_872_sll_83 <= 0;
      __delay_data_876__variable_76 <= 0;
      __delay_data_880_eq_95 <= 0;
      __delay_data_873__delay_872_sll_83 <= 0;
      __delay_data_877__delay_876__variable_76 <= 0;
      __delay_data_881__delay_880_eq_95 <= 0;
      __delay_data_874__delay_873__delay_872_sll_83 <= 0;
      __delay_data_878__delay_877__delay_876__variable_76 <= 0;
      __delay_data_882__delay_881__delay_880_eq_95 <= 0;
      __delay_data_875__delay_874__delay_873__delay_872_sll_83 <= 0;
      __delay_data_879__delay_878__delay_877__delay_876__variable_76 <= 0;
      __delay_data_883__delay_882__delay_881__delay_880_eq_95 <= 0;
      _cond_data_96 <= 0;
      _greaterthan_data_97 <= 0;
      _lessthan_data_101 <= 0;
      _greatereq_data_105 <= 0;
      __delay_data_884_cond_96 <= 0;
      _cond_data_99 <= 0;
      _cond_data_103 <= 0;
      __delay_data_885_greatereq_105 <= 0;
      _cond_data_107 <= 0;
      __variable_wdata_74 <= 0;
      __variable_wdata_75 <= 0;
      __variable_wdata_76 <= 0;
      _tmp_1122 <= 0;
      _tmp_1123 <= 0;
      _tmp_1124 <= 0;
      _tmp_1125 <= 0;
      _tmp_1126 <= 0;
      _tmp_1127 <= 0;
      _tmp_1128 <= 0;
      _tmp_1129 <= 0;
      _tmp_1130 <= 0;
      _tmp_1131 <= 0;
      _tmp_1132 <= 0;
      _tmp_1133 <= 0;
      _tmp_1134 <= 0;
      _tmp_1135 <= 0;
      _tmp_1136 <= 0;
      _tmp_1137 <= 0;
      _tmp_1138 <= 0;
      _tmp_1139 <= 0;
      _tmp_1140 <= 0;
      _tmp_1141 <= 0;
      _tmp_1142 <= 0;
      _tmp_1143 <= 0;
      _tmp_1144 <= 0;
      _tmp_1145 <= 0;
      _tmp_1146 <= 0;
      _tmp_1147 <= 0;
      _tmp_1148 <= 0;
      _tmp_1149 <= 0;
      _tmp_1150 <= 0;
      _tmp_1151 <= 0;
      _tmp_1152 <= 0;
      _tmp_1153 <= 0;
      _tmp_1154 <= 0;
      _tmp_1155 <= 0;
      _mul_rshift_round_clip_4_busy_reg <= 0;
    end else begin
      if(_mul_rshift_round_clip_4_stream_oready) begin
        _mul_rshift_round_clip_4_x_source_ram_renable <= 0;
        _mul_rshift_round_clip_4_x_source_fifo_deq <= 0;
      end 
      _mul_rshift_round_clip_4_x_idle <= _mul_rshift_round_clip_4_x_idle;
      if(_mul_rshift_round_clip_4_stream_oready) begin
        _mul_rshift_round_clip_4_y_source_ram_renable <= 0;
        _mul_rshift_round_clip_4_y_source_fifo_deq <= 0;
      end 
      _mul_rshift_round_clip_4_y_idle <= _mul_rshift_round_clip_4_y_idle;
      if(_mul_rshift_round_clip_4_stream_oready) begin
        _mul_rshift_round_clip_4_rshift_source_ram_renable <= 0;
        _mul_rshift_round_clip_4_rshift_source_fifo_deq <= 0;
      end 
      _mul_rshift_round_clip_4_rshift_idle <= _mul_rshift_round_clip_4_rshift_idle;
      if(_mul_rshift_round_clip_4_stream_oready) begin
        _mul_rshift_round_clip_4_z_sink_wenable <= 0;
        _mul_rshift_round_clip_4_z_sink_fifo_enq <= 0;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        __mul_rshift_round_clip_4_stream_ivalid_1 <= _mul_rshift_round_clip_4_stream_ivalid;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        __mul_rshift_round_clip_4_stream_ivalid_2 <= __mul_rshift_round_clip_4_stream_ivalid_1;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        __mul_rshift_round_clip_4_stream_ivalid_3 <= __mul_rshift_round_clip_4_stream_ivalid_2;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        __mul_rshift_round_clip_4_stream_ivalid_4 <= __mul_rshift_round_clip_4_stream_ivalid_3;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        __mul_rshift_round_clip_4_stream_ivalid_5 <= __mul_rshift_round_clip_4_stream_ivalid_4;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        __mul_rshift_round_clip_4_stream_ivalid_6 <= __mul_rshift_round_clip_4_stream_ivalid_5;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        __mul_rshift_round_clip_4_stream_ivalid_7 <= __mul_rshift_round_clip_4_stream_ivalid_6;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        __mul_rshift_round_clip_4_stream_ivalid_8 <= __mul_rshift_round_clip_4_stream_ivalid_7;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        _times_mul_odata_reg_77 <= _times_mul_odata_77;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        __delay_data_872_sll_83 <= _sll_data_83;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        __delay_data_876__variable_76 <= mul_rshift_round_clip_4_rshift_data;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        __delay_data_880_eq_95 <= _eq_data_95;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        __delay_data_873__delay_872_sll_83 <= __delay_data_872_sll_83;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        __delay_data_877__delay_876__variable_76 <= __delay_data_876__variable_76;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        __delay_data_881__delay_880_eq_95 <= __delay_data_880_eq_95;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        __delay_data_874__delay_873__delay_872_sll_83 <= __delay_data_873__delay_872_sll_83;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        __delay_data_878__delay_877__delay_876__variable_76 <= __delay_data_877__delay_876__variable_76;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        __delay_data_882__delay_881__delay_880_eq_95 <= __delay_data_881__delay_880_eq_95;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        __delay_data_875__delay_874__delay_873__delay_872_sll_83 <= __delay_data_874__delay_873__delay_872_sll_83;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        __delay_data_879__delay_878__delay_877__delay_876__variable_76 <= __delay_data_878__delay_877__delay_876__variable_76;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        __delay_data_883__delay_882__delay_881__delay_880_eq_95 <= __delay_data_882__delay_881__delay_880_eq_95;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        _cond_data_96 <= (__delay_data_883__delay_882__delay_881__delay_880_eq_95)? _times_data_77 : _sra_data_93;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        _greaterthan_data_97 <= _cond_data_96 > 8'sd127;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        _lessthan_data_101 <= _cond_data_96 < -8'sd127;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        _greatereq_data_105 <= _cond_data_96 >= 1'sd0;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        __delay_data_884_cond_96 <= _cond_data_96;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        _cond_data_99 <= (_greaterthan_data_97)? 8'sd127 : __delay_data_884_cond_96;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        _cond_data_103 <= (_lessthan_data_101)? -8'sd127 : __delay_data_884_cond_96;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        __delay_data_885_greatereq_105 <= _greatereq_data_105;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        _cond_data_107 <= (__delay_data_885_greatereq_105)? _cond_data_99 : _cond_data_103;
      end 
      if(__stream_conv2d_24_stream_ivalid_20 && _stream_conv2d_24_stream_oready) begin
        __variable_wdata_74 <= _plus_data_870;
      end 
      if(__stream_conv2d_24_stream_ivalid_20 && _stream_conv2d_24_stream_oready) begin
        __variable_wdata_75 <= __delay_data_1141__delay_1140__delay_1139__delay_1138___cond_332;
      end 
      if(__stream_conv2d_24_stream_ivalid_20 && _stream_conv2d_24_stream_oready) begin
        __variable_wdata_76 <= __delay_data_1160__delay_1159__delay_1158__delay_1157___plus_886;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        _tmp_1122 <= _mul_rshift_round_clip_4_source_start;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        _tmp_1123 <= _tmp_1122;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        _tmp_1124 <= _tmp_1123;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        _tmp_1125 <= _mul_rshift_round_clip_4_source_start;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        _tmp_1126 <= _tmp_1125;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        _tmp_1127 <= _tmp_1126;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        _tmp_1128 <= _tmp_1127;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        _tmp_1129 <= _tmp_1128;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        _tmp_1130 <= _tmp_1129;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        _tmp_1131 <= _tmp_1130;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        _tmp_1132 <= _tmp_1131;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        _tmp_1133 <= _tmp_1132;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        _tmp_1134 <= _tmp_1133;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        _tmp_1135 <= _mul_rshift_round_clip_4_source_stop;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        _tmp_1136 <= _tmp_1135;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        _tmp_1137 <= _tmp_1136;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        _tmp_1138 <= _tmp_1137;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        _tmp_1139 <= _tmp_1138;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        _tmp_1140 <= _tmp_1139;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        _tmp_1141 <= _tmp_1140;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        _tmp_1142 <= _tmp_1141;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        _tmp_1143 <= _tmp_1142;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        _tmp_1144 <= _tmp_1143;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        _tmp_1145 <= _mul_rshift_round_clip_4_source_busy;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        _tmp_1146 <= _tmp_1145;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        _tmp_1147 <= _tmp_1146;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        _tmp_1148 <= _tmp_1147;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        _tmp_1149 <= _tmp_1148;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        _tmp_1150 <= _tmp_1149;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        _tmp_1151 <= _tmp_1150;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        _tmp_1152 <= _tmp_1151;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        _tmp_1153 <= _tmp_1152;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        _tmp_1154 <= _tmp_1153;
      end 
      if(_mul_rshift_round_clip_4_stream_oready) begin
        _tmp_1155 <= _mul_rshift_round_clip_4_sink_busy;
      end 
      if(!_mul_rshift_round_clip_4_sink_busy && _tmp_1155) begin
        _mul_rshift_round_clip_4_busy_reg <= 0;
      end 
      if(_mul_rshift_round_clip_4_source_busy) begin
        _mul_rshift_round_clip_4_busy_reg <= 1;
      end 
      if(__stream_matmul_55_stream_ivalid_18 && _stream_matmul_55_stream_oready) begin
        __variable_wdata_74 <= _plus_data_1023;
      end 
      if(__stream_matmul_55_stream_ivalid_18 && _stream_matmul_55_stream_oready) begin
        __variable_wdata_75 <= __delay_data_1261__delay_1260__delay_1259__delay_1258___cond_964;
      end 
      if(__stream_matmul_55_stream_ivalid_18 && _stream_matmul_55_stream_oready) begin
        __variable_wdata_76 <= __delay_data_1278__delay_1277__delay_1276___plus_1025;
      end 
    end
  end

  localparam _mul_rshift_round_clip_4_fsm_1 = 1;
  localparam _mul_rshift_round_clip_4_fsm_2 = 2;
  localparam _mul_rshift_round_clip_4_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_rshift_round_clip_4_fsm <= _mul_rshift_round_clip_4_fsm_init;
      _mul_rshift_round_clip_4_source_start <= 0;
      _mul_rshift_round_clip_4_source_busy <= 0;
      _mul_rshift_round_clip_4_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_24_stream_ivalid_20 && _stream_conv2d_24_stream_oready) begin
        _mul_rshift_round_clip_4_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_24_stream_oready && _stream_conv2d_24_busy) begin
        _mul_rshift_round_clip_4_source_busy <= _stream_conv2d_24_source_busy;
      end 
      if(_mul_rshift_round_clip_4_stream_oready && _tmp_1124) begin
        _mul_rshift_round_clip_4_stream_ivalid <= 1;
      end 
      if(_mul_rshift_round_clip_4_stream_oready && 1'd0) begin
        _mul_rshift_round_clip_4_stream_ivalid <= 0;
      end 
      if(__stream_matmul_55_stream_ivalid_18 && _stream_matmul_55_stream_oready) begin
        _mul_rshift_round_clip_4_stream_ivalid <= 1'd1;
      end 
      if(_stream_matmul_55_stream_oready && _stream_matmul_55_busy) begin
        _mul_rshift_round_clip_4_source_busy <= _stream_matmul_55_source_busy;
      end 
      case(_mul_rshift_round_clip_4_fsm)
        _mul_rshift_round_clip_4_fsm_init: begin
          if(_mul_rshift_round_clip_4_run_flag) begin
            _mul_rshift_round_clip_4_source_start <= 1;
          end 
          if(_mul_rshift_round_clip_4_run_flag) begin
            _mul_rshift_round_clip_4_fsm <= _mul_rshift_round_clip_4_fsm_1;
          end 
        end
        _mul_rshift_round_clip_4_fsm_1: begin
          if(_mul_rshift_round_clip_4_source_start && _mul_rshift_round_clip_4_stream_oready) begin
            _mul_rshift_round_clip_4_source_start <= 0;
            _mul_rshift_round_clip_4_source_busy <= 1;
          end 
          if(_mul_rshift_round_clip_4_source_start && _mul_rshift_round_clip_4_stream_oready) begin
            _mul_rshift_round_clip_4_fsm <= _mul_rshift_round_clip_4_fsm_2;
          end 
        end
        _mul_rshift_round_clip_4_fsm_2: begin
          if(_mul_rshift_round_clip_4_stream_oready) begin
            _mul_rshift_round_clip_4_fsm <= _mul_rshift_round_clip_4_fsm_3;
          end 
        end
        _mul_rshift_round_clip_4_fsm_3: begin
          if(_mul_rshift_round_clip_4_stream_oready && 1'd0) begin
            _mul_rshift_round_clip_4_source_busy <= 0;
          end 
          if(_mul_rshift_round_clip_4_stream_oready && 1'd0 && _mul_rshift_round_clip_4_run_flag) begin
            _mul_rshift_round_clip_4_source_start <= 1;
          end 
          if(_mul_rshift_round_clip_4_stream_oready && 1'd0) begin
            _mul_rshift_round_clip_4_fsm <= _mul_rshift_round_clip_4_fsm_init;
          end 
          if(_mul_rshift_round_clip_4_stream_oready && 1'd0 && _mul_rshift_round_clip_4_run_flag) begin
            _mul_rshift_round_clip_4_fsm <= _mul_rshift_round_clip_4_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_5_x_source_ram_renable <= 0;
      _mul_5_x_source_fifo_deq <= 0;
      _mul_5_x_idle <= 1;
      _mul_5_y_source_ram_renable <= 0;
      _mul_5_y_source_fifo_deq <= 0;
      _mul_5_y_idle <= 1;
      _mul_5_rshift_source_ram_renable <= 0;
      _mul_5_rshift_source_fifo_deq <= 0;
      _mul_5_rshift_idle <= 1;
      _mul_5_z_sink_wenable <= 0;
      _mul_5_z_sink_fifo_enq <= 0;
      __mul_5_stream_ivalid_1 <= 0;
      __mul_5_stream_ivalid_2 <= 0;
      __mul_5_stream_ivalid_3 <= 0;
      __mul_5_stream_ivalid_4 <= 0;
      __mul_5_stream_ivalid_5 <= 0;
      __mul_5_stream_ivalid_6 <= 0;
      __mul_5_stream_ivalid_7 <= 0;
      __mul_5_stream_ivalid_8 <= 0;
      _greaterthan_data_111 <= 0;
      _minus_data_113 <= 0;
      _greatereq_data_124 <= 0;
      __delay_data_686__variable_108 <= 0;
      __delay_data_689__variable_109 <= 0;
      __delay_data_692__variable_110 <= 0;
      _sll_data_115 <= 0;
      __delay_data_683_greaterthan_111 <= 0;
      __delay_data_684_greatereq_124 <= 0;
      __delay_data_687__delay_686__variable_108 <= 0;
      __delay_data_690__delay_689__variable_109 <= 0;
      __delay_data_693__delay_692__variable_110 <= 0;
      _cond_data_121 <= 0;
      __delay_data_685__delay_684_greatereq_124 <= 0;
      __delay_data_688__delay_687__delay_686__variable_108 <= 0;
      __delay_data_691__delay_690__delay_689__variable_109 <= 0;
      __delay_data_694__delay_693__delay_692__variable_110 <= 0;
      __muladd_madd_odata_reg_127 <= 0;
      __delay_data_695__delay_694__delay_693____variable_110 <= 0;
      __delay_data_696__delay_695__delay_694____variable_110 <= 0;
      __delay_data_697__delay_696__delay_695____variable_110 <= 0;
      __delay_data_698__delay_697__delay_696____variable_110 <= 0;
      _sra_data_128 <= 0;
      __variable_wdata_108 <= 0;
      __variable_wdata_109 <= 0;
      __variable_wdata_110 <= 0;
      _tmp_768 <= 0;
      _tmp_769 <= 0;
      _tmp_770 <= 0;
      _tmp_771 <= 0;
      _tmp_772 <= 0;
      _tmp_773 <= 0;
      _tmp_774 <= 0;
      _tmp_775 <= 0;
      _tmp_776 <= 0;
      _tmp_777 <= 0;
      _tmp_778 <= 0;
      _tmp_779 <= 0;
      _tmp_780 <= 0;
      _tmp_781 <= 0;
      _tmp_782 <= 0;
      _tmp_783 <= 0;
      _tmp_784 <= 0;
      _tmp_785 <= 0;
      _tmp_786 <= 0;
      _tmp_787 <= 0;
      _tmp_788 <= 0;
      _tmp_789 <= 0;
      _tmp_790 <= 0;
      _tmp_791 <= 0;
      _tmp_792 <= 0;
      _tmp_793 <= 0;
      _tmp_794 <= 0;
      _tmp_795 <= 0;
      _tmp_796 <= 0;
      _tmp_797 <= 0;
      _tmp_798 <= 0;
      _tmp_799 <= 0;
      _tmp_800 <= 0;
      _tmp_801 <= 0;
      _mul_5_busy_reg <= 0;
    end else begin
      if(_mul_5_stream_oready) begin
        _mul_5_x_source_ram_renable <= 0;
        _mul_5_x_source_fifo_deq <= 0;
      end 
      _mul_5_x_idle <= _mul_5_x_idle;
      if(_mul_5_stream_oready) begin
        _mul_5_y_source_ram_renable <= 0;
        _mul_5_y_source_fifo_deq <= 0;
      end 
      _mul_5_y_idle <= _mul_5_y_idle;
      if(_mul_5_stream_oready) begin
        _mul_5_rshift_source_ram_renable <= 0;
        _mul_5_rshift_source_fifo_deq <= 0;
      end 
      _mul_5_rshift_idle <= _mul_5_rshift_idle;
      if(_mul_5_stream_oready) begin
        _mul_5_z_sink_wenable <= 0;
        _mul_5_z_sink_fifo_enq <= 0;
      end 
      if(_mul_5_stream_oready) begin
        __mul_5_stream_ivalid_1 <= _mul_5_stream_ivalid;
      end 
      if(_mul_5_stream_oready) begin
        __mul_5_stream_ivalid_2 <= __mul_5_stream_ivalid_1;
      end 
      if(_mul_5_stream_oready) begin
        __mul_5_stream_ivalid_3 <= __mul_5_stream_ivalid_2;
      end 
      if(_mul_5_stream_oready) begin
        __mul_5_stream_ivalid_4 <= __mul_5_stream_ivalid_3;
      end 
      if(_mul_5_stream_oready) begin
        __mul_5_stream_ivalid_5 <= __mul_5_stream_ivalid_4;
      end 
      if(_mul_5_stream_oready) begin
        __mul_5_stream_ivalid_6 <= __mul_5_stream_ivalid_5;
      end 
      if(_mul_5_stream_oready) begin
        __mul_5_stream_ivalid_7 <= __mul_5_stream_ivalid_6;
      end 
      if(_mul_5_stream_oready) begin
        __mul_5_stream_ivalid_8 <= __mul_5_stream_ivalid_7;
      end 
      if(_mul_5_stream_oready) begin
        _greaterthan_data_111 <= mul_5_rshift_data > 1'sd0;
      end 
      if(_mul_5_stream_oready) begin
        _minus_data_113 <= mul_5_rshift_data - 2'sd1;
      end 
      if(_mul_5_stream_oready) begin
        _greatereq_data_124 <= mul_5_x_data >= 1'sd0;
      end 
      if(_mul_5_stream_oready) begin
        __delay_data_686__variable_108 <= mul_5_x_data;
      end 
      if(_mul_5_stream_oready) begin
        __delay_data_689__variable_109 <= mul_5_y_data;
      end 
      if(_mul_5_stream_oready) begin
        __delay_data_692__variable_110 <= mul_5_rshift_data;
      end 
      if(_mul_5_stream_oready) begin
        _sll_data_115 <= 2'sd1 << _minus_data_113;
      end 
      if(_mul_5_stream_oready) begin
        __delay_data_683_greaterthan_111 <= _greaterthan_data_111;
      end 
      if(_mul_5_stream_oready) begin
        __delay_data_684_greatereq_124 <= _greatereq_data_124;
      end 
      if(_mul_5_stream_oready) begin
        __delay_data_687__delay_686__variable_108 <= __delay_data_686__variable_108;
      end 
      if(_mul_5_stream_oready) begin
        __delay_data_690__delay_689__variable_109 <= __delay_data_689__variable_109;
      end 
      if(_mul_5_stream_oready) begin
        __delay_data_693__delay_692__variable_110 <= __delay_data_692__variable_110;
      end 
      if(_mul_5_stream_oready) begin
        _cond_data_121 <= (__delay_data_683_greaterthan_111)? _sll_data_115 : 1'sd0;
      end 
      if(_mul_5_stream_oready) begin
        __delay_data_685__delay_684_greatereq_124 <= __delay_data_684_greatereq_124;
      end 
      if(_mul_5_stream_oready) begin
        __delay_data_688__delay_687__delay_686__variable_108 <= __delay_data_687__delay_686__variable_108;
      end 
      if(_mul_5_stream_oready) begin
        __delay_data_691__delay_690__delay_689__variable_109 <= __delay_data_690__delay_689__variable_109;
      end 
      if(_mul_5_stream_oready) begin
        __delay_data_694__delay_693__delay_692__variable_110 <= __delay_data_693__delay_692__variable_110;
      end 
      if(_mul_5_stream_oready) begin
        __muladd_madd_odata_reg_127 <= __muladd_madd_odata_127;
      end 
      if(_mul_5_stream_oready) begin
        __delay_data_695__delay_694__delay_693____variable_110 <= __delay_data_694__delay_693__delay_692__variable_110;
      end 
      if(_mul_5_stream_oready) begin
        __delay_data_696__delay_695__delay_694____variable_110 <= __delay_data_695__delay_694__delay_693____variable_110;
      end 
      if(_mul_5_stream_oready) begin
        __delay_data_697__delay_696__delay_695____variable_110 <= __delay_data_696__delay_695__delay_694____variable_110;
      end 
      if(_mul_5_stream_oready) begin
        __delay_data_698__delay_697__delay_696____variable_110 <= __delay_data_697__delay_696__delay_695____variable_110;
      end 
      if(_mul_5_stream_oready) begin
        _sra_data_128 <= __muladd_data_127 >>> __delay_data_698__delay_697__delay_696____variable_110;
      end 
      if(__stream_conv2d_24_stream_ivalid_1 && _stream_conv2d_24_stream_oready) begin
        __variable_wdata_108 <= _cond_data_665;
      end 
      if(__stream_conv2d_24_stream_ivalid_1 && _stream_conv2d_24_stream_oready) begin
        __variable_wdata_109 <= __delay_data_1048_reinterpretcast_637;
      end 
      if(__stream_conv2d_24_stream_ivalid_1 && _stream_conv2d_24_stream_oready) begin
        __variable_wdata_110 <= _plus_data_699;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_768 <= _mul_5_source_start;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_769 <= _tmp_768;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_770 <= _tmp_769;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_771 <= _mul_5_source_start;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_772 <= _tmp_771;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_773 <= _tmp_772;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_774 <= _tmp_773;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_775 <= _tmp_774;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_776 <= _tmp_775;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_777 <= _tmp_776;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_778 <= _tmp_777;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_779 <= _tmp_778;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_780 <= _tmp_779;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_781 <= _mul_5_source_stop;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_782 <= _tmp_781;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_783 <= _tmp_782;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_784 <= _tmp_783;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_785 <= _tmp_784;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_786 <= _tmp_785;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_787 <= _tmp_786;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_788 <= _tmp_787;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_789 <= _tmp_788;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_790 <= _tmp_789;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_791 <= _mul_5_source_busy;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_792 <= _tmp_791;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_793 <= _tmp_792;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_794 <= _tmp_793;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_795 <= _tmp_794;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_796 <= _tmp_795;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_797 <= _tmp_796;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_798 <= _tmp_797;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_799 <= _tmp_798;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_800 <= _tmp_799;
      end 
      if(_mul_5_stream_oready) begin
        _tmp_801 <= _mul_5_sink_busy;
      end 
      if(!_mul_5_sink_busy && _tmp_801) begin
        _mul_5_busy_reg <= 0;
      end 
      if(_mul_5_source_busy) begin
        _mul_5_busy_reg <= 1;
      end 
      if(__stream_matmul_55_stream_ivalid_1 && _stream_matmul_55_stream_oready) begin
        __variable_wdata_108 <= _cond_data_1013;
      end 
      if(__stream_matmul_55_stream_ivalid_1 && _stream_matmul_55_stream_oready) begin
        __variable_wdata_109 <= __delay_data_1194_reinterpretcast_1009;
      end 
      if(__stream_matmul_55_stream_ivalid_1 && _stream_matmul_55_stream_oready) begin
        __variable_wdata_110 <= _plus_data_1015;
      end 
    end
  end

  localparam _mul_5_fsm_1 = 1;
  localparam _mul_5_fsm_2 = 2;
  localparam _mul_5_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_5_fsm <= _mul_5_fsm_init;
      _mul_5_source_start <= 0;
      _mul_5_source_busy <= 0;
      _mul_5_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_24_stream_ivalid_1 && _stream_conv2d_24_stream_oready) begin
        _mul_5_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_24_stream_oready && _stream_conv2d_24_busy) begin
        _mul_5_source_busy <= _stream_conv2d_24_source_busy;
      end 
      if(_mul_5_stream_oready && _tmp_770) begin
        _mul_5_stream_ivalid <= 1;
      end 
      if(_mul_5_stream_oready && 1'd0) begin
        _mul_5_stream_ivalid <= 0;
      end 
      if(__stream_matmul_55_stream_ivalid_1 && _stream_matmul_55_stream_oready) begin
        _mul_5_stream_ivalid <= 1'd1;
      end 
      if(_stream_matmul_55_stream_oready && _stream_matmul_55_busy) begin
        _mul_5_source_busy <= _stream_matmul_55_source_busy;
      end 
      case(_mul_5_fsm)
        _mul_5_fsm_init: begin
          if(_mul_5_run_flag) begin
            _mul_5_source_start <= 1;
          end 
          if(_mul_5_run_flag) begin
            _mul_5_fsm <= _mul_5_fsm_1;
          end 
        end
        _mul_5_fsm_1: begin
          if(_mul_5_source_start && _mul_5_stream_oready) begin
            _mul_5_source_start <= 0;
            _mul_5_source_busy <= 1;
          end 
          if(_mul_5_source_start && _mul_5_stream_oready) begin
            _mul_5_fsm <= _mul_5_fsm_2;
          end 
        end
        _mul_5_fsm_2: begin
          if(_mul_5_stream_oready) begin
            _mul_5_fsm <= _mul_5_fsm_3;
          end 
        end
        _mul_5_fsm_3: begin
          if(_mul_5_stream_oready && 1'd0) begin
            _mul_5_source_busy <= 0;
          end 
          if(_mul_5_stream_oready && 1'd0 && _mul_5_run_flag) begin
            _mul_5_source_start <= 1;
          end 
          if(_mul_5_stream_oready && 1'd0) begin
            _mul_5_fsm <= _mul_5_fsm_init;
          end 
          if(_mul_5_stream_oready && 1'd0 && _mul_5_run_flag) begin
            _mul_5_fsm <= _mul_5_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_6_x_source_ram_renable <= 0;
      _mul_6_x_source_fifo_deq <= 0;
      _mul_6_x_idle <= 1;
      _mul_6_y_source_ram_renable <= 0;
      _mul_6_y_source_fifo_deq <= 0;
      _mul_6_y_idle <= 1;
      _mul_6_rshift_source_ram_renable <= 0;
      _mul_6_rshift_source_fifo_deq <= 0;
      _mul_6_rshift_idle <= 1;
      _mul_6_z_sink_wenable <= 0;
      _mul_6_z_sink_fifo_enq <= 0;
      __mul_6_stream_ivalid_1 <= 0;
      __mul_6_stream_ivalid_2 <= 0;
      __mul_6_stream_ivalid_3 <= 0;
      __mul_6_stream_ivalid_4 <= 0;
      __mul_6_stream_ivalid_5 <= 0;
      __mul_6_stream_ivalid_6 <= 0;
      __mul_6_stream_ivalid_7 <= 0;
      __mul_6_stream_ivalid_8 <= 0;
      _greaterthan_data_132 <= 0;
      _minus_data_134 <= 0;
      _greatereq_data_145 <= 0;
      __delay_data_705__variable_129 <= 0;
      __delay_data_708__variable_130 <= 0;
      __delay_data_711__variable_131 <= 0;
      _sll_data_136 <= 0;
      __delay_data_702_greaterthan_132 <= 0;
      __delay_data_703_greatereq_145 <= 0;
      __delay_data_706__delay_705__variable_129 <= 0;
      __delay_data_709__delay_708__variable_130 <= 0;
      __delay_data_712__delay_711__variable_131 <= 0;
      _cond_data_142 <= 0;
      __delay_data_704__delay_703_greatereq_145 <= 0;
      __delay_data_707__delay_706__delay_705__variable_129 <= 0;
      __delay_data_710__delay_709__delay_708__variable_130 <= 0;
      __delay_data_713__delay_712__delay_711__variable_131 <= 0;
      __muladd_madd_odata_reg_148 <= 0;
      __delay_data_714__delay_713__delay_712____variable_131 <= 0;
      __delay_data_715__delay_714__delay_713____variable_131 <= 0;
      __delay_data_716__delay_715__delay_714____variable_131 <= 0;
      __delay_data_717__delay_716__delay_715____variable_131 <= 0;
      _sra_data_149 <= 0;
      __variable_wdata_129 <= 0;
      __variable_wdata_130 <= 0;
      __variable_wdata_131 <= 0;
      _tmp_802 <= 0;
      _tmp_803 <= 0;
      _tmp_804 <= 0;
      _tmp_805 <= 0;
      _tmp_806 <= 0;
      _tmp_807 <= 0;
      _tmp_808 <= 0;
      _tmp_809 <= 0;
      _tmp_810 <= 0;
      _tmp_811 <= 0;
      _tmp_812 <= 0;
      _tmp_813 <= 0;
      _tmp_814 <= 0;
      _tmp_815 <= 0;
      _tmp_816 <= 0;
      _tmp_817 <= 0;
      _tmp_818 <= 0;
      _tmp_819 <= 0;
      _tmp_820 <= 0;
      _tmp_821 <= 0;
      _tmp_822 <= 0;
      _tmp_823 <= 0;
      _tmp_824 <= 0;
      _tmp_825 <= 0;
      _tmp_826 <= 0;
      _tmp_827 <= 0;
      _tmp_828 <= 0;
      _tmp_829 <= 0;
      _tmp_830 <= 0;
      _tmp_831 <= 0;
      _tmp_832 <= 0;
      _tmp_833 <= 0;
      _tmp_834 <= 0;
      _tmp_835 <= 0;
      _mul_6_busy_reg <= 0;
    end else begin
      if(_mul_6_stream_oready) begin
        _mul_6_x_source_ram_renable <= 0;
        _mul_6_x_source_fifo_deq <= 0;
      end 
      _mul_6_x_idle <= _mul_6_x_idle;
      if(_mul_6_stream_oready) begin
        _mul_6_y_source_ram_renable <= 0;
        _mul_6_y_source_fifo_deq <= 0;
      end 
      _mul_6_y_idle <= _mul_6_y_idle;
      if(_mul_6_stream_oready) begin
        _mul_6_rshift_source_ram_renable <= 0;
        _mul_6_rshift_source_fifo_deq <= 0;
      end 
      _mul_6_rshift_idle <= _mul_6_rshift_idle;
      if(_mul_6_stream_oready) begin
        _mul_6_z_sink_wenable <= 0;
        _mul_6_z_sink_fifo_enq <= 0;
      end 
      if(_mul_6_stream_oready) begin
        __mul_6_stream_ivalid_1 <= _mul_6_stream_ivalid;
      end 
      if(_mul_6_stream_oready) begin
        __mul_6_stream_ivalid_2 <= __mul_6_stream_ivalid_1;
      end 
      if(_mul_6_stream_oready) begin
        __mul_6_stream_ivalid_3 <= __mul_6_stream_ivalid_2;
      end 
      if(_mul_6_stream_oready) begin
        __mul_6_stream_ivalid_4 <= __mul_6_stream_ivalid_3;
      end 
      if(_mul_6_stream_oready) begin
        __mul_6_stream_ivalid_5 <= __mul_6_stream_ivalid_4;
      end 
      if(_mul_6_stream_oready) begin
        __mul_6_stream_ivalid_6 <= __mul_6_stream_ivalid_5;
      end 
      if(_mul_6_stream_oready) begin
        __mul_6_stream_ivalid_7 <= __mul_6_stream_ivalid_6;
      end 
      if(_mul_6_stream_oready) begin
        __mul_6_stream_ivalid_8 <= __mul_6_stream_ivalid_7;
      end 
      if(_mul_6_stream_oready) begin
        _greaterthan_data_132 <= mul_6_rshift_data > 1'sd0;
      end 
      if(_mul_6_stream_oready) begin
        _minus_data_134 <= mul_6_rshift_data - 2'sd1;
      end 
      if(_mul_6_stream_oready) begin
        _greatereq_data_145 <= mul_6_x_data >= 1'sd0;
      end 
      if(_mul_6_stream_oready) begin
        __delay_data_705__variable_129 <= mul_6_x_data;
      end 
      if(_mul_6_stream_oready) begin
        __delay_data_708__variable_130 <= mul_6_y_data;
      end 
      if(_mul_6_stream_oready) begin
        __delay_data_711__variable_131 <= mul_6_rshift_data;
      end 
      if(_mul_6_stream_oready) begin
        _sll_data_136 <= 2'sd1 << _minus_data_134;
      end 
      if(_mul_6_stream_oready) begin
        __delay_data_702_greaterthan_132 <= _greaterthan_data_132;
      end 
      if(_mul_6_stream_oready) begin
        __delay_data_703_greatereq_145 <= _greatereq_data_145;
      end 
      if(_mul_6_stream_oready) begin
        __delay_data_706__delay_705__variable_129 <= __delay_data_705__variable_129;
      end 
      if(_mul_6_stream_oready) begin
        __delay_data_709__delay_708__variable_130 <= __delay_data_708__variable_130;
      end 
      if(_mul_6_stream_oready) begin
        __delay_data_712__delay_711__variable_131 <= __delay_data_711__variable_131;
      end 
      if(_mul_6_stream_oready) begin
        _cond_data_142 <= (__delay_data_702_greaterthan_132)? _sll_data_136 : 1'sd0;
      end 
      if(_mul_6_stream_oready) begin
        __delay_data_704__delay_703_greatereq_145 <= __delay_data_703_greatereq_145;
      end 
      if(_mul_6_stream_oready) begin
        __delay_data_707__delay_706__delay_705__variable_129 <= __delay_data_706__delay_705__variable_129;
      end 
      if(_mul_6_stream_oready) begin
        __delay_data_710__delay_709__delay_708__variable_130 <= __delay_data_709__delay_708__variable_130;
      end 
      if(_mul_6_stream_oready) begin
        __delay_data_713__delay_712__delay_711__variable_131 <= __delay_data_712__delay_711__variable_131;
      end 
      if(_mul_6_stream_oready) begin
        __muladd_madd_odata_reg_148 <= __muladd_madd_odata_148;
      end 
      if(_mul_6_stream_oready) begin
        __delay_data_714__delay_713__delay_712____variable_131 <= __delay_data_713__delay_712__delay_711__variable_131;
      end 
      if(_mul_6_stream_oready) begin
        __delay_data_715__delay_714__delay_713____variable_131 <= __delay_data_714__delay_713__delay_712____variable_131;
      end 
      if(_mul_6_stream_oready) begin
        __delay_data_716__delay_715__delay_714____variable_131 <= __delay_data_715__delay_714__delay_713____variable_131;
      end 
      if(_mul_6_stream_oready) begin
        __delay_data_717__delay_716__delay_715____variable_131 <= __delay_data_716__delay_715__delay_714____variable_131;
      end 
      if(_mul_6_stream_oready) begin
        _sra_data_149 <= __muladd_data_148 >>> __delay_data_717__delay_716__delay_715____variable_131;
      end 
      if(__stream_conv2d_24_stream_ivalid_1 && _stream_conv2d_24_stream_oready) begin
        __variable_wdata_129 <= _cond_data_667;
      end 
      if(__stream_conv2d_24_stream_ivalid_1 && _stream_conv2d_24_stream_oready) begin
        __variable_wdata_130 <= __delay_data_1050_reinterpretcast_638;
      end 
      if(__stream_conv2d_24_stream_ivalid_1 && _stream_conv2d_24_stream_oready) begin
        __variable_wdata_131 <= _plus_data_718;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_802 <= _mul_6_source_start;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_803 <= _tmp_802;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_804 <= _tmp_803;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_805 <= _mul_6_source_start;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_806 <= _tmp_805;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_807 <= _tmp_806;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_808 <= _tmp_807;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_809 <= _tmp_808;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_810 <= _tmp_809;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_811 <= _tmp_810;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_812 <= _tmp_811;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_813 <= _tmp_812;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_814 <= _tmp_813;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_815 <= _mul_6_source_stop;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_816 <= _tmp_815;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_817 <= _tmp_816;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_818 <= _tmp_817;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_819 <= _tmp_818;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_820 <= _tmp_819;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_821 <= _tmp_820;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_822 <= _tmp_821;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_823 <= _tmp_822;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_824 <= _tmp_823;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_825 <= _mul_6_source_busy;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_826 <= _tmp_825;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_827 <= _tmp_826;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_828 <= _tmp_827;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_829 <= _tmp_828;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_830 <= _tmp_829;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_831 <= _tmp_830;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_832 <= _tmp_831;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_833 <= _tmp_832;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_834 <= _tmp_833;
      end 
      if(_mul_6_stream_oready) begin
        _tmp_835 <= _mul_6_sink_busy;
      end 
      if(!_mul_6_sink_busy && _tmp_835) begin
        _mul_6_busy_reg <= 0;
      end 
      if(_mul_6_source_busy) begin
        _mul_6_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_6_fsm_1 = 1;
  localparam _mul_6_fsm_2 = 2;
  localparam _mul_6_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_6_fsm <= _mul_6_fsm_init;
      _mul_6_source_start <= 0;
      _mul_6_source_busy <= 0;
      _mul_6_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_24_stream_ivalid_1 && _stream_conv2d_24_stream_oready) begin
        _mul_6_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_24_stream_oready && _stream_conv2d_24_busy) begin
        _mul_6_source_busy <= _stream_conv2d_24_source_busy;
      end 
      if(_mul_6_stream_oready && _tmp_804) begin
        _mul_6_stream_ivalid <= 1;
      end 
      if(_mul_6_stream_oready && 1'd0) begin
        _mul_6_stream_ivalid <= 0;
      end 
      case(_mul_6_fsm)
        _mul_6_fsm_init: begin
          if(_mul_6_run_flag) begin
            _mul_6_source_start <= 1;
          end 
          if(_mul_6_run_flag) begin
            _mul_6_fsm <= _mul_6_fsm_1;
          end 
        end
        _mul_6_fsm_1: begin
          if(_mul_6_source_start && _mul_6_stream_oready) begin
            _mul_6_source_start <= 0;
            _mul_6_source_busy <= 1;
          end 
          if(_mul_6_source_start && _mul_6_stream_oready) begin
            _mul_6_fsm <= _mul_6_fsm_2;
          end 
        end
        _mul_6_fsm_2: begin
          if(_mul_6_stream_oready) begin
            _mul_6_fsm <= _mul_6_fsm_3;
          end 
        end
        _mul_6_fsm_3: begin
          if(_mul_6_stream_oready && 1'd0) begin
            _mul_6_source_busy <= 0;
          end 
          if(_mul_6_stream_oready && 1'd0 && _mul_6_run_flag) begin
            _mul_6_source_start <= 1;
          end 
          if(_mul_6_stream_oready && 1'd0) begin
            _mul_6_fsm <= _mul_6_fsm_init;
          end 
          if(_mul_6_stream_oready && 1'd0 && _mul_6_run_flag) begin
            _mul_6_fsm <= _mul_6_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_7_x_source_ram_renable <= 0;
      _mul_7_x_source_fifo_deq <= 0;
      _mul_7_x_idle <= 1;
      _mul_7_y_source_ram_renable <= 0;
      _mul_7_y_source_fifo_deq <= 0;
      _mul_7_y_idle <= 1;
      _mul_7_rshift_source_ram_renable <= 0;
      _mul_7_rshift_source_fifo_deq <= 0;
      _mul_7_rshift_idle <= 1;
      _mul_7_z_sink_wenable <= 0;
      _mul_7_z_sink_fifo_enq <= 0;
      __mul_7_stream_ivalid_1 <= 0;
      __mul_7_stream_ivalid_2 <= 0;
      __mul_7_stream_ivalid_3 <= 0;
      __mul_7_stream_ivalid_4 <= 0;
      __mul_7_stream_ivalid_5 <= 0;
      __mul_7_stream_ivalid_6 <= 0;
      __mul_7_stream_ivalid_7 <= 0;
      __mul_7_stream_ivalid_8 <= 0;
      _greaterthan_data_153 <= 0;
      _minus_data_155 <= 0;
      _greatereq_data_166 <= 0;
      __delay_data_724__variable_150 <= 0;
      __delay_data_727__variable_151 <= 0;
      __delay_data_730__variable_152 <= 0;
      _sll_data_157 <= 0;
      __delay_data_721_greaterthan_153 <= 0;
      __delay_data_722_greatereq_166 <= 0;
      __delay_data_725__delay_724__variable_150 <= 0;
      __delay_data_728__delay_727__variable_151 <= 0;
      __delay_data_731__delay_730__variable_152 <= 0;
      _cond_data_163 <= 0;
      __delay_data_723__delay_722_greatereq_166 <= 0;
      __delay_data_726__delay_725__delay_724__variable_150 <= 0;
      __delay_data_729__delay_728__delay_727__variable_151 <= 0;
      __delay_data_732__delay_731__delay_730__variable_152 <= 0;
      __muladd_madd_odata_reg_169 <= 0;
      __delay_data_733__delay_732__delay_731____variable_152 <= 0;
      __delay_data_734__delay_733__delay_732____variable_152 <= 0;
      __delay_data_735__delay_734__delay_733____variable_152 <= 0;
      __delay_data_736__delay_735__delay_734____variable_152 <= 0;
      _sra_data_170 <= 0;
      __variable_wdata_150 <= 0;
      __variable_wdata_151 <= 0;
      __variable_wdata_152 <= 0;
      _tmp_836 <= 0;
      _tmp_837 <= 0;
      _tmp_838 <= 0;
      _tmp_839 <= 0;
      _tmp_840 <= 0;
      _tmp_841 <= 0;
      _tmp_842 <= 0;
      _tmp_843 <= 0;
      _tmp_844 <= 0;
      _tmp_845 <= 0;
      _tmp_846 <= 0;
      _tmp_847 <= 0;
      _tmp_848 <= 0;
      _tmp_849 <= 0;
      _tmp_850 <= 0;
      _tmp_851 <= 0;
      _tmp_852 <= 0;
      _tmp_853 <= 0;
      _tmp_854 <= 0;
      _tmp_855 <= 0;
      _tmp_856 <= 0;
      _tmp_857 <= 0;
      _tmp_858 <= 0;
      _tmp_859 <= 0;
      _tmp_860 <= 0;
      _tmp_861 <= 0;
      _tmp_862 <= 0;
      _tmp_863 <= 0;
      _tmp_864 <= 0;
      _tmp_865 <= 0;
      _tmp_866 <= 0;
      _tmp_867 <= 0;
      _tmp_868 <= 0;
      _tmp_869 <= 0;
      _mul_7_busy_reg <= 0;
    end else begin
      if(_mul_7_stream_oready) begin
        _mul_7_x_source_ram_renable <= 0;
        _mul_7_x_source_fifo_deq <= 0;
      end 
      _mul_7_x_idle <= _mul_7_x_idle;
      if(_mul_7_stream_oready) begin
        _mul_7_y_source_ram_renable <= 0;
        _mul_7_y_source_fifo_deq <= 0;
      end 
      _mul_7_y_idle <= _mul_7_y_idle;
      if(_mul_7_stream_oready) begin
        _mul_7_rshift_source_ram_renable <= 0;
        _mul_7_rshift_source_fifo_deq <= 0;
      end 
      _mul_7_rshift_idle <= _mul_7_rshift_idle;
      if(_mul_7_stream_oready) begin
        _mul_7_z_sink_wenable <= 0;
        _mul_7_z_sink_fifo_enq <= 0;
      end 
      if(_mul_7_stream_oready) begin
        __mul_7_stream_ivalid_1 <= _mul_7_stream_ivalid;
      end 
      if(_mul_7_stream_oready) begin
        __mul_7_stream_ivalid_2 <= __mul_7_stream_ivalid_1;
      end 
      if(_mul_7_stream_oready) begin
        __mul_7_stream_ivalid_3 <= __mul_7_stream_ivalid_2;
      end 
      if(_mul_7_stream_oready) begin
        __mul_7_stream_ivalid_4 <= __mul_7_stream_ivalid_3;
      end 
      if(_mul_7_stream_oready) begin
        __mul_7_stream_ivalid_5 <= __mul_7_stream_ivalid_4;
      end 
      if(_mul_7_stream_oready) begin
        __mul_7_stream_ivalid_6 <= __mul_7_stream_ivalid_5;
      end 
      if(_mul_7_stream_oready) begin
        __mul_7_stream_ivalid_7 <= __mul_7_stream_ivalid_6;
      end 
      if(_mul_7_stream_oready) begin
        __mul_7_stream_ivalid_8 <= __mul_7_stream_ivalid_7;
      end 
      if(_mul_7_stream_oready) begin
        _greaterthan_data_153 <= mul_7_rshift_data > 1'sd0;
      end 
      if(_mul_7_stream_oready) begin
        _minus_data_155 <= mul_7_rshift_data - 2'sd1;
      end 
      if(_mul_7_stream_oready) begin
        _greatereq_data_166 <= mul_7_x_data >= 1'sd0;
      end 
      if(_mul_7_stream_oready) begin
        __delay_data_724__variable_150 <= mul_7_x_data;
      end 
      if(_mul_7_stream_oready) begin
        __delay_data_727__variable_151 <= mul_7_y_data;
      end 
      if(_mul_7_stream_oready) begin
        __delay_data_730__variable_152 <= mul_7_rshift_data;
      end 
      if(_mul_7_stream_oready) begin
        _sll_data_157 <= 2'sd1 << _minus_data_155;
      end 
      if(_mul_7_stream_oready) begin
        __delay_data_721_greaterthan_153 <= _greaterthan_data_153;
      end 
      if(_mul_7_stream_oready) begin
        __delay_data_722_greatereq_166 <= _greatereq_data_166;
      end 
      if(_mul_7_stream_oready) begin
        __delay_data_725__delay_724__variable_150 <= __delay_data_724__variable_150;
      end 
      if(_mul_7_stream_oready) begin
        __delay_data_728__delay_727__variable_151 <= __delay_data_727__variable_151;
      end 
      if(_mul_7_stream_oready) begin
        __delay_data_731__delay_730__variable_152 <= __delay_data_730__variable_152;
      end 
      if(_mul_7_stream_oready) begin
        _cond_data_163 <= (__delay_data_721_greaterthan_153)? _sll_data_157 : 1'sd0;
      end 
      if(_mul_7_stream_oready) begin
        __delay_data_723__delay_722_greatereq_166 <= __delay_data_722_greatereq_166;
      end 
      if(_mul_7_stream_oready) begin
        __delay_data_726__delay_725__delay_724__variable_150 <= __delay_data_725__delay_724__variable_150;
      end 
      if(_mul_7_stream_oready) begin
        __delay_data_729__delay_728__delay_727__variable_151 <= __delay_data_728__delay_727__variable_151;
      end 
      if(_mul_7_stream_oready) begin
        __delay_data_732__delay_731__delay_730__variable_152 <= __delay_data_731__delay_730__variable_152;
      end 
      if(_mul_7_stream_oready) begin
        __muladd_madd_odata_reg_169 <= __muladd_madd_odata_169;
      end 
      if(_mul_7_stream_oready) begin
        __delay_data_733__delay_732__delay_731____variable_152 <= __delay_data_732__delay_731__delay_730__variable_152;
      end 
      if(_mul_7_stream_oready) begin
        __delay_data_734__delay_733__delay_732____variable_152 <= __delay_data_733__delay_732__delay_731____variable_152;
      end 
      if(_mul_7_stream_oready) begin
        __delay_data_735__delay_734__delay_733____variable_152 <= __delay_data_734__delay_733__delay_732____variable_152;
      end 
      if(_mul_7_stream_oready) begin
        __delay_data_736__delay_735__delay_734____variable_152 <= __delay_data_735__delay_734__delay_733____variable_152;
      end 
      if(_mul_7_stream_oready) begin
        _sra_data_170 <= __muladd_data_169 >>> __delay_data_736__delay_735__delay_734____variable_152;
      end 
      if(__stream_conv2d_24_stream_ivalid_1 && _stream_conv2d_24_stream_oready) begin
        __variable_wdata_150 <= _cond_data_669;
      end 
      if(__stream_conv2d_24_stream_ivalid_1 && _stream_conv2d_24_stream_oready) begin
        __variable_wdata_151 <= __delay_data_1052_reinterpretcast_639;
      end 
      if(__stream_conv2d_24_stream_ivalid_1 && _stream_conv2d_24_stream_oready) begin
        __variable_wdata_152 <= _plus_data_737;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_836 <= _mul_7_source_start;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_837 <= _tmp_836;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_838 <= _tmp_837;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_839 <= _mul_7_source_start;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_840 <= _tmp_839;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_841 <= _tmp_840;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_842 <= _tmp_841;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_843 <= _tmp_842;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_844 <= _tmp_843;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_845 <= _tmp_844;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_846 <= _tmp_845;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_847 <= _tmp_846;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_848 <= _tmp_847;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_849 <= _mul_7_source_stop;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_850 <= _tmp_849;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_851 <= _tmp_850;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_852 <= _tmp_851;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_853 <= _tmp_852;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_854 <= _tmp_853;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_855 <= _tmp_854;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_856 <= _tmp_855;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_857 <= _tmp_856;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_858 <= _tmp_857;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_859 <= _mul_7_source_busy;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_860 <= _tmp_859;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_861 <= _tmp_860;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_862 <= _tmp_861;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_863 <= _tmp_862;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_864 <= _tmp_863;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_865 <= _tmp_864;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_866 <= _tmp_865;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_867 <= _tmp_866;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_868 <= _tmp_867;
      end 
      if(_mul_7_stream_oready) begin
        _tmp_869 <= _mul_7_sink_busy;
      end 
      if(!_mul_7_sink_busy && _tmp_869) begin
        _mul_7_busy_reg <= 0;
      end 
      if(_mul_7_source_busy) begin
        _mul_7_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_7_fsm_1 = 1;
  localparam _mul_7_fsm_2 = 2;
  localparam _mul_7_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_7_fsm <= _mul_7_fsm_init;
      _mul_7_source_start <= 0;
      _mul_7_source_busy <= 0;
      _mul_7_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_24_stream_ivalid_1 && _stream_conv2d_24_stream_oready) begin
        _mul_7_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_24_stream_oready && _stream_conv2d_24_busy) begin
        _mul_7_source_busy <= _stream_conv2d_24_source_busy;
      end 
      if(_mul_7_stream_oready && _tmp_838) begin
        _mul_7_stream_ivalid <= 1;
      end 
      if(_mul_7_stream_oready && 1'd0) begin
        _mul_7_stream_ivalid <= 0;
      end 
      case(_mul_7_fsm)
        _mul_7_fsm_init: begin
          if(_mul_7_run_flag) begin
            _mul_7_source_start <= 1;
          end 
          if(_mul_7_run_flag) begin
            _mul_7_fsm <= _mul_7_fsm_1;
          end 
        end
        _mul_7_fsm_1: begin
          if(_mul_7_source_start && _mul_7_stream_oready) begin
            _mul_7_source_start <= 0;
            _mul_7_source_busy <= 1;
          end 
          if(_mul_7_source_start && _mul_7_stream_oready) begin
            _mul_7_fsm <= _mul_7_fsm_2;
          end 
        end
        _mul_7_fsm_2: begin
          if(_mul_7_stream_oready) begin
            _mul_7_fsm <= _mul_7_fsm_3;
          end 
        end
        _mul_7_fsm_3: begin
          if(_mul_7_stream_oready && 1'd0) begin
            _mul_7_source_busy <= 0;
          end 
          if(_mul_7_stream_oready && 1'd0 && _mul_7_run_flag) begin
            _mul_7_source_start <= 1;
          end 
          if(_mul_7_stream_oready && 1'd0) begin
            _mul_7_fsm <= _mul_7_fsm_init;
          end 
          if(_mul_7_stream_oready && 1'd0 && _mul_7_run_flag) begin
            _mul_7_fsm <= _mul_7_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_8_x_source_ram_renable <= 0;
      _mul_8_x_source_fifo_deq <= 0;
      _mul_8_x_idle <= 1;
      _mul_8_y_source_ram_renable <= 0;
      _mul_8_y_source_fifo_deq <= 0;
      _mul_8_y_idle <= 1;
      _mul_8_rshift_source_ram_renable <= 0;
      _mul_8_rshift_source_fifo_deq <= 0;
      _mul_8_rshift_idle <= 1;
      _mul_8_z_sink_wenable <= 0;
      _mul_8_z_sink_fifo_enq <= 0;
      __mul_8_stream_ivalid_1 <= 0;
      __mul_8_stream_ivalid_2 <= 0;
      __mul_8_stream_ivalid_3 <= 0;
      __mul_8_stream_ivalid_4 <= 0;
      __mul_8_stream_ivalid_5 <= 0;
      __mul_8_stream_ivalid_6 <= 0;
      __mul_8_stream_ivalid_7 <= 0;
      __mul_8_stream_ivalid_8 <= 0;
      _greaterthan_data_174 <= 0;
      _minus_data_176 <= 0;
      _greatereq_data_187 <= 0;
      __delay_data_743__variable_171 <= 0;
      __delay_data_746__variable_172 <= 0;
      __delay_data_749__variable_173 <= 0;
      _sll_data_178 <= 0;
      __delay_data_740_greaterthan_174 <= 0;
      __delay_data_741_greatereq_187 <= 0;
      __delay_data_744__delay_743__variable_171 <= 0;
      __delay_data_747__delay_746__variable_172 <= 0;
      __delay_data_750__delay_749__variable_173 <= 0;
      _cond_data_184 <= 0;
      __delay_data_742__delay_741_greatereq_187 <= 0;
      __delay_data_745__delay_744__delay_743__variable_171 <= 0;
      __delay_data_748__delay_747__delay_746__variable_172 <= 0;
      __delay_data_751__delay_750__delay_749__variable_173 <= 0;
      __muladd_madd_odata_reg_190 <= 0;
      __delay_data_752__delay_751__delay_750____variable_173 <= 0;
      __delay_data_753__delay_752__delay_751____variable_173 <= 0;
      __delay_data_754__delay_753__delay_752____variable_173 <= 0;
      __delay_data_755__delay_754__delay_753____variable_173 <= 0;
      _sra_data_191 <= 0;
      __variable_wdata_171 <= 0;
      __variable_wdata_172 <= 0;
      __variable_wdata_173 <= 0;
      _tmp_870 <= 0;
      _tmp_871 <= 0;
      _tmp_872 <= 0;
      _tmp_873 <= 0;
      _tmp_874 <= 0;
      _tmp_875 <= 0;
      _tmp_876 <= 0;
      _tmp_877 <= 0;
      _tmp_878 <= 0;
      _tmp_879 <= 0;
      _tmp_880 <= 0;
      _tmp_881 <= 0;
      _tmp_882 <= 0;
      _tmp_883 <= 0;
      _tmp_884 <= 0;
      _tmp_885 <= 0;
      _tmp_886 <= 0;
      _tmp_887 <= 0;
      _tmp_888 <= 0;
      _tmp_889 <= 0;
      _tmp_890 <= 0;
      _tmp_891 <= 0;
      _tmp_892 <= 0;
      _tmp_893 <= 0;
      _tmp_894 <= 0;
      _tmp_895 <= 0;
      _tmp_896 <= 0;
      _tmp_897 <= 0;
      _tmp_898 <= 0;
      _tmp_899 <= 0;
      _tmp_900 <= 0;
      _tmp_901 <= 0;
      _tmp_902 <= 0;
      _tmp_903 <= 0;
      _mul_8_busy_reg <= 0;
    end else begin
      if(_mul_8_stream_oready) begin
        _mul_8_x_source_ram_renable <= 0;
        _mul_8_x_source_fifo_deq <= 0;
      end 
      _mul_8_x_idle <= _mul_8_x_idle;
      if(_mul_8_stream_oready) begin
        _mul_8_y_source_ram_renable <= 0;
        _mul_8_y_source_fifo_deq <= 0;
      end 
      _mul_8_y_idle <= _mul_8_y_idle;
      if(_mul_8_stream_oready) begin
        _mul_8_rshift_source_ram_renable <= 0;
        _mul_8_rshift_source_fifo_deq <= 0;
      end 
      _mul_8_rshift_idle <= _mul_8_rshift_idle;
      if(_mul_8_stream_oready) begin
        _mul_8_z_sink_wenable <= 0;
        _mul_8_z_sink_fifo_enq <= 0;
      end 
      if(_mul_8_stream_oready) begin
        __mul_8_stream_ivalid_1 <= _mul_8_stream_ivalid;
      end 
      if(_mul_8_stream_oready) begin
        __mul_8_stream_ivalid_2 <= __mul_8_stream_ivalid_1;
      end 
      if(_mul_8_stream_oready) begin
        __mul_8_stream_ivalid_3 <= __mul_8_stream_ivalid_2;
      end 
      if(_mul_8_stream_oready) begin
        __mul_8_stream_ivalid_4 <= __mul_8_stream_ivalid_3;
      end 
      if(_mul_8_stream_oready) begin
        __mul_8_stream_ivalid_5 <= __mul_8_stream_ivalid_4;
      end 
      if(_mul_8_stream_oready) begin
        __mul_8_stream_ivalid_6 <= __mul_8_stream_ivalid_5;
      end 
      if(_mul_8_stream_oready) begin
        __mul_8_stream_ivalid_7 <= __mul_8_stream_ivalid_6;
      end 
      if(_mul_8_stream_oready) begin
        __mul_8_stream_ivalid_8 <= __mul_8_stream_ivalid_7;
      end 
      if(_mul_8_stream_oready) begin
        _greaterthan_data_174 <= mul_8_rshift_data > 1'sd0;
      end 
      if(_mul_8_stream_oready) begin
        _minus_data_176 <= mul_8_rshift_data - 2'sd1;
      end 
      if(_mul_8_stream_oready) begin
        _greatereq_data_187 <= mul_8_x_data >= 1'sd0;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_743__variable_171 <= mul_8_x_data;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_746__variable_172 <= mul_8_y_data;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_749__variable_173 <= mul_8_rshift_data;
      end 
      if(_mul_8_stream_oready) begin
        _sll_data_178 <= 2'sd1 << _minus_data_176;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_740_greaterthan_174 <= _greaterthan_data_174;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_741_greatereq_187 <= _greatereq_data_187;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_744__delay_743__variable_171 <= __delay_data_743__variable_171;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_747__delay_746__variable_172 <= __delay_data_746__variable_172;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_750__delay_749__variable_173 <= __delay_data_749__variable_173;
      end 
      if(_mul_8_stream_oready) begin
        _cond_data_184 <= (__delay_data_740_greaterthan_174)? _sll_data_178 : 1'sd0;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_742__delay_741_greatereq_187 <= __delay_data_741_greatereq_187;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_745__delay_744__delay_743__variable_171 <= __delay_data_744__delay_743__variable_171;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_748__delay_747__delay_746__variable_172 <= __delay_data_747__delay_746__variable_172;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_751__delay_750__delay_749__variable_173 <= __delay_data_750__delay_749__variable_173;
      end 
      if(_mul_8_stream_oready) begin
        __muladd_madd_odata_reg_190 <= __muladd_madd_odata_190;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_752__delay_751__delay_750____variable_173 <= __delay_data_751__delay_750__delay_749__variable_173;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_753__delay_752__delay_751____variable_173 <= __delay_data_752__delay_751__delay_750____variable_173;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_754__delay_753__delay_752____variable_173 <= __delay_data_753__delay_752__delay_751____variable_173;
      end 
      if(_mul_8_stream_oready) begin
        __delay_data_755__delay_754__delay_753____variable_173 <= __delay_data_754__delay_753__delay_752____variable_173;
      end 
      if(_mul_8_stream_oready) begin
        _sra_data_191 <= __muladd_data_190 >>> __delay_data_755__delay_754__delay_753____variable_173;
      end 
      if(__stream_conv2d_24_stream_ivalid_1 && _stream_conv2d_24_stream_oready) begin
        __variable_wdata_171 <= _cond_data_671;
      end 
      if(__stream_conv2d_24_stream_ivalid_1 && _stream_conv2d_24_stream_oready) begin
        __variable_wdata_172 <= __delay_data_1054_reinterpretcast_640;
      end 
      if(__stream_conv2d_24_stream_ivalid_1 && _stream_conv2d_24_stream_oready) begin
        __variable_wdata_173 <= _plus_data_756;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_870 <= _mul_8_source_start;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_871 <= _tmp_870;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_872 <= _tmp_871;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_873 <= _mul_8_source_start;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_874 <= _tmp_873;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_875 <= _tmp_874;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_876 <= _tmp_875;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_877 <= _tmp_876;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_878 <= _tmp_877;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_879 <= _tmp_878;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_880 <= _tmp_879;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_881 <= _tmp_880;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_882 <= _tmp_881;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_883 <= _mul_8_source_stop;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_884 <= _tmp_883;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_885 <= _tmp_884;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_886 <= _tmp_885;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_887 <= _tmp_886;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_888 <= _tmp_887;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_889 <= _tmp_888;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_890 <= _tmp_889;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_891 <= _tmp_890;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_892 <= _tmp_891;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_893 <= _mul_8_source_busy;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_894 <= _tmp_893;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_895 <= _tmp_894;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_896 <= _tmp_895;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_897 <= _tmp_896;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_898 <= _tmp_897;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_899 <= _tmp_898;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_900 <= _tmp_899;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_901 <= _tmp_900;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_902 <= _tmp_901;
      end 
      if(_mul_8_stream_oready) begin
        _tmp_903 <= _mul_8_sink_busy;
      end 
      if(!_mul_8_sink_busy && _tmp_903) begin
        _mul_8_busy_reg <= 0;
      end 
      if(_mul_8_source_busy) begin
        _mul_8_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_8_fsm_1 = 1;
  localparam _mul_8_fsm_2 = 2;
  localparam _mul_8_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_8_fsm <= _mul_8_fsm_init;
      _mul_8_source_start <= 0;
      _mul_8_source_busy <= 0;
      _mul_8_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_24_stream_ivalid_1 && _stream_conv2d_24_stream_oready) begin
        _mul_8_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_24_stream_oready && _stream_conv2d_24_busy) begin
        _mul_8_source_busy <= _stream_conv2d_24_source_busy;
      end 
      if(_mul_8_stream_oready && _tmp_872) begin
        _mul_8_stream_ivalid <= 1;
      end 
      if(_mul_8_stream_oready && 1'd0) begin
        _mul_8_stream_ivalid <= 0;
      end 
      case(_mul_8_fsm)
        _mul_8_fsm_init: begin
          if(_mul_8_run_flag) begin
            _mul_8_source_start <= 1;
          end 
          if(_mul_8_run_flag) begin
            _mul_8_fsm <= _mul_8_fsm_1;
          end 
        end
        _mul_8_fsm_1: begin
          if(_mul_8_source_start && _mul_8_stream_oready) begin
            _mul_8_source_start <= 0;
            _mul_8_source_busy <= 1;
          end 
          if(_mul_8_source_start && _mul_8_stream_oready) begin
            _mul_8_fsm <= _mul_8_fsm_2;
          end 
        end
        _mul_8_fsm_2: begin
          if(_mul_8_stream_oready) begin
            _mul_8_fsm <= _mul_8_fsm_3;
          end 
        end
        _mul_8_fsm_3: begin
          if(_mul_8_stream_oready && 1'd0) begin
            _mul_8_source_busy <= 0;
          end 
          if(_mul_8_stream_oready && 1'd0 && _mul_8_run_flag) begin
            _mul_8_source_start <= 1;
          end 
          if(_mul_8_stream_oready && 1'd0) begin
            _mul_8_fsm <= _mul_8_fsm_init;
          end 
          if(_mul_8_stream_oready && 1'd0 && _mul_8_run_flag) begin
            _mul_8_fsm <= _mul_8_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_9_x_source_ram_renable <= 0;
      _mul_9_x_source_fifo_deq <= 0;
      _mul_9_x_idle <= 1;
      _mul_9_y_source_ram_renable <= 0;
      _mul_9_y_source_fifo_deq <= 0;
      _mul_9_y_idle <= 1;
      _mul_9_rshift_source_ram_renable <= 0;
      _mul_9_rshift_source_fifo_deq <= 0;
      _mul_9_rshift_idle <= 1;
      _mul_9_z_sink_wenable <= 0;
      _mul_9_z_sink_fifo_enq <= 0;
      __mul_9_stream_ivalid_1 <= 0;
      __mul_9_stream_ivalid_2 <= 0;
      __mul_9_stream_ivalid_3 <= 0;
      __mul_9_stream_ivalid_4 <= 0;
      __mul_9_stream_ivalid_5 <= 0;
      __mul_9_stream_ivalid_6 <= 0;
      __mul_9_stream_ivalid_7 <= 0;
      __mul_9_stream_ivalid_8 <= 0;
      _greaterthan_data_195 <= 0;
      _minus_data_197 <= 0;
      _greatereq_data_208 <= 0;
      __delay_data_762__variable_192 <= 0;
      __delay_data_765__variable_193 <= 0;
      __delay_data_768__variable_194 <= 0;
      _sll_data_199 <= 0;
      __delay_data_759_greaterthan_195 <= 0;
      __delay_data_760_greatereq_208 <= 0;
      __delay_data_763__delay_762__variable_192 <= 0;
      __delay_data_766__delay_765__variable_193 <= 0;
      __delay_data_769__delay_768__variable_194 <= 0;
      _cond_data_205 <= 0;
      __delay_data_761__delay_760_greatereq_208 <= 0;
      __delay_data_764__delay_763__delay_762__variable_192 <= 0;
      __delay_data_767__delay_766__delay_765__variable_193 <= 0;
      __delay_data_770__delay_769__delay_768__variable_194 <= 0;
      __muladd_madd_odata_reg_211 <= 0;
      __delay_data_771__delay_770__delay_769____variable_194 <= 0;
      __delay_data_772__delay_771__delay_770____variable_194 <= 0;
      __delay_data_773__delay_772__delay_771____variable_194 <= 0;
      __delay_data_774__delay_773__delay_772____variable_194 <= 0;
      _sra_data_212 <= 0;
      __variable_wdata_192 <= 0;
      __variable_wdata_193 <= 0;
      __variable_wdata_194 <= 0;
      _tmp_904 <= 0;
      _tmp_905 <= 0;
      _tmp_906 <= 0;
      _tmp_907 <= 0;
      _tmp_908 <= 0;
      _tmp_909 <= 0;
      _tmp_910 <= 0;
      _tmp_911 <= 0;
      _tmp_912 <= 0;
      _tmp_913 <= 0;
      _tmp_914 <= 0;
      _tmp_915 <= 0;
      _tmp_916 <= 0;
      _tmp_917 <= 0;
      _tmp_918 <= 0;
      _tmp_919 <= 0;
      _tmp_920 <= 0;
      _tmp_921 <= 0;
      _tmp_922 <= 0;
      _tmp_923 <= 0;
      _tmp_924 <= 0;
      _tmp_925 <= 0;
      _tmp_926 <= 0;
      _tmp_927 <= 0;
      _tmp_928 <= 0;
      _tmp_929 <= 0;
      _tmp_930 <= 0;
      _tmp_931 <= 0;
      _tmp_932 <= 0;
      _tmp_933 <= 0;
      _tmp_934 <= 0;
      _tmp_935 <= 0;
      _tmp_936 <= 0;
      _tmp_937 <= 0;
      _mul_9_busy_reg <= 0;
    end else begin
      if(_mul_9_stream_oready) begin
        _mul_9_x_source_ram_renable <= 0;
        _mul_9_x_source_fifo_deq <= 0;
      end 
      _mul_9_x_idle <= _mul_9_x_idle;
      if(_mul_9_stream_oready) begin
        _mul_9_y_source_ram_renable <= 0;
        _mul_9_y_source_fifo_deq <= 0;
      end 
      _mul_9_y_idle <= _mul_9_y_idle;
      if(_mul_9_stream_oready) begin
        _mul_9_rshift_source_ram_renable <= 0;
        _mul_9_rshift_source_fifo_deq <= 0;
      end 
      _mul_9_rshift_idle <= _mul_9_rshift_idle;
      if(_mul_9_stream_oready) begin
        _mul_9_z_sink_wenable <= 0;
        _mul_9_z_sink_fifo_enq <= 0;
      end 
      if(_mul_9_stream_oready) begin
        __mul_9_stream_ivalid_1 <= _mul_9_stream_ivalid;
      end 
      if(_mul_9_stream_oready) begin
        __mul_9_stream_ivalid_2 <= __mul_9_stream_ivalid_1;
      end 
      if(_mul_9_stream_oready) begin
        __mul_9_stream_ivalid_3 <= __mul_9_stream_ivalid_2;
      end 
      if(_mul_9_stream_oready) begin
        __mul_9_stream_ivalid_4 <= __mul_9_stream_ivalid_3;
      end 
      if(_mul_9_stream_oready) begin
        __mul_9_stream_ivalid_5 <= __mul_9_stream_ivalid_4;
      end 
      if(_mul_9_stream_oready) begin
        __mul_9_stream_ivalid_6 <= __mul_9_stream_ivalid_5;
      end 
      if(_mul_9_stream_oready) begin
        __mul_9_stream_ivalid_7 <= __mul_9_stream_ivalid_6;
      end 
      if(_mul_9_stream_oready) begin
        __mul_9_stream_ivalid_8 <= __mul_9_stream_ivalid_7;
      end 
      if(_mul_9_stream_oready) begin
        _greaterthan_data_195 <= mul_9_rshift_data > 1'sd0;
      end 
      if(_mul_9_stream_oready) begin
        _minus_data_197 <= mul_9_rshift_data - 2'sd1;
      end 
      if(_mul_9_stream_oready) begin
        _greatereq_data_208 <= mul_9_x_data >= 1'sd0;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_762__variable_192 <= mul_9_x_data;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_765__variable_193 <= mul_9_y_data;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_768__variable_194 <= mul_9_rshift_data;
      end 
      if(_mul_9_stream_oready) begin
        _sll_data_199 <= 2'sd1 << _minus_data_197;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_759_greaterthan_195 <= _greaterthan_data_195;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_760_greatereq_208 <= _greatereq_data_208;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_763__delay_762__variable_192 <= __delay_data_762__variable_192;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_766__delay_765__variable_193 <= __delay_data_765__variable_193;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_769__delay_768__variable_194 <= __delay_data_768__variable_194;
      end 
      if(_mul_9_stream_oready) begin
        _cond_data_205 <= (__delay_data_759_greaterthan_195)? _sll_data_199 : 1'sd0;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_761__delay_760_greatereq_208 <= __delay_data_760_greatereq_208;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_764__delay_763__delay_762__variable_192 <= __delay_data_763__delay_762__variable_192;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_767__delay_766__delay_765__variable_193 <= __delay_data_766__delay_765__variable_193;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_770__delay_769__delay_768__variable_194 <= __delay_data_769__delay_768__variable_194;
      end 
      if(_mul_9_stream_oready) begin
        __muladd_madd_odata_reg_211 <= __muladd_madd_odata_211;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_771__delay_770__delay_769____variable_194 <= __delay_data_770__delay_769__delay_768__variable_194;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_772__delay_771__delay_770____variable_194 <= __delay_data_771__delay_770__delay_769____variable_194;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_773__delay_772__delay_771____variable_194 <= __delay_data_772__delay_771__delay_770____variable_194;
      end 
      if(_mul_9_stream_oready) begin
        __delay_data_774__delay_773__delay_772____variable_194 <= __delay_data_773__delay_772__delay_771____variable_194;
      end 
      if(_mul_9_stream_oready) begin
        _sra_data_212 <= __muladd_data_211 >>> __delay_data_774__delay_773__delay_772____variable_194;
      end 
      if(__stream_conv2d_24_stream_ivalid_1 && _stream_conv2d_24_stream_oready) begin
        __variable_wdata_192 <= _cond_data_673;
      end 
      if(__stream_conv2d_24_stream_ivalid_1 && _stream_conv2d_24_stream_oready) begin
        __variable_wdata_193 <= __delay_data_1056_reinterpretcast_641;
      end 
      if(__stream_conv2d_24_stream_ivalid_1 && _stream_conv2d_24_stream_oready) begin
        __variable_wdata_194 <= _plus_data_775;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_904 <= _mul_9_source_start;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_905 <= _tmp_904;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_906 <= _tmp_905;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_907 <= _mul_9_source_start;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_908 <= _tmp_907;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_909 <= _tmp_908;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_910 <= _tmp_909;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_911 <= _tmp_910;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_912 <= _tmp_911;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_913 <= _tmp_912;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_914 <= _tmp_913;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_915 <= _tmp_914;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_916 <= _tmp_915;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_917 <= _mul_9_source_stop;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_918 <= _tmp_917;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_919 <= _tmp_918;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_920 <= _tmp_919;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_921 <= _tmp_920;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_922 <= _tmp_921;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_923 <= _tmp_922;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_924 <= _tmp_923;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_925 <= _tmp_924;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_926 <= _tmp_925;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_927 <= _mul_9_source_busy;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_928 <= _tmp_927;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_929 <= _tmp_928;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_930 <= _tmp_929;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_931 <= _tmp_930;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_932 <= _tmp_931;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_933 <= _tmp_932;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_934 <= _tmp_933;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_935 <= _tmp_934;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_936 <= _tmp_935;
      end 
      if(_mul_9_stream_oready) begin
        _tmp_937 <= _mul_9_sink_busy;
      end 
      if(!_mul_9_sink_busy && _tmp_937) begin
        _mul_9_busy_reg <= 0;
      end 
      if(_mul_9_source_busy) begin
        _mul_9_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_9_fsm_1 = 1;
  localparam _mul_9_fsm_2 = 2;
  localparam _mul_9_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_9_fsm <= _mul_9_fsm_init;
      _mul_9_source_start <= 0;
      _mul_9_source_busy <= 0;
      _mul_9_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_24_stream_ivalid_1 && _stream_conv2d_24_stream_oready) begin
        _mul_9_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_24_stream_oready && _stream_conv2d_24_busy) begin
        _mul_9_source_busy <= _stream_conv2d_24_source_busy;
      end 
      if(_mul_9_stream_oready && _tmp_906) begin
        _mul_9_stream_ivalid <= 1;
      end 
      if(_mul_9_stream_oready && 1'd0) begin
        _mul_9_stream_ivalid <= 0;
      end 
      case(_mul_9_fsm)
        _mul_9_fsm_init: begin
          if(_mul_9_run_flag) begin
            _mul_9_source_start <= 1;
          end 
          if(_mul_9_run_flag) begin
            _mul_9_fsm <= _mul_9_fsm_1;
          end 
        end
        _mul_9_fsm_1: begin
          if(_mul_9_source_start && _mul_9_stream_oready) begin
            _mul_9_source_start <= 0;
            _mul_9_source_busy <= 1;
          end 
          if(_mul_9_source_start && _mul_9_stream_oready) begin
            _mul_9_fsm <= _mul_9_fsm_2;
          end 
        end
        _mul_9_fsm_2: begin
          if(_mul_9_stream_oready) begin
            _mul_9_fsm <= _mul_9_fsm_3;
          end 
        end
        _mul_9_fsm_3: begin
          if(_mul_9_stream_oready && 1'd0) begin
            _mul_9_source_busy <= 0;
          end 
          if(_mul_9_stream_oready && 1'd0 && _mul_9_run_flag) begin
            _mul_9_source_start <= 1;
          end 
          if(_mul_9_stream_oready && 1'd0) begin
            _mul_9_fsm <= _mul_9_fsm_init;
          end 
          if(_mul_9_stream_oready && 1'd0 && _mul_9_run_flag) begin
            _mul_9_fsm <= _mul_9_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_10_x_source_ram_renable <= 0;
      _mul_10_x_source_fifo_deq <= 0;
      _mul_10_x_idle <= 1;
      _mul_10_y_source_ram_renable <= 0;
      _mul_10_y_source_fifo_deq <= 0;
      _mul_10_y_idle <= 1;
      _mul_10_rshift_source_ram_renable <= 0;
      _mul_10_rshift_source_fifo_deq <= 0;
      _mul_10_rshift_idle <= 1;
      _mul_10_z_sink_wenable <= 0;
      _mul_10_z_sink_fifo_enq <= 0;
      __mul_10_stream_ivalid_1 <= 0;
      __mul_10_stream_ivalid_2 <= 0;
      __mul_10_stream_ivalid_3 <= 0;
      __mul_10_stream_ivalid_4 <= 0;
      __mul_10_stream_ivalid_5 <= 0;
      __mul_10_stream_ivalid_6 <= 0;
      __mul_10_stream_ivalid_7 <= 0;
      __mul_10_stream_ivalid_8 <= 0;
      _greaterthan_data_216 <= 0;
      _minus_data_218 <= 0;
      _greatereq_data_229 <= 0;
      __delay_data_781__variable_213 <= 0;
      __delay_data_784__variable_214 <= 0;
      __delay_data_787__variable_215 <= 0;
      _sll_data_220 <= 0;
      __delay_data_778_greaterthan_216 <= 0;
      __delay_data_779_greatereq_229 <= 0;
      __delay_data_782__delay_781__variable_213 <= 0;
      __delay_data_785__delay_784__variable_214 <= 0;
      __delay_data_788__delay_787__variable_215 <= 0;
      _cond_data_226 <= 0;
      __delay_data_780__delay_779_greatereq_229 <= 0;
      __delay_data_783__delay_782__delay_781__variable_213 <= 0;
      __delay_data_786__delay_785__delay_784__variable_214 <= 0;
      __delay_data_789__delay_788__delay_787__variable_215 <= 0;
      __muladd_madd_odata_reg_232 <= 0;
      __delay_data_790__delay_789__delay_788____variable_215 <= 0;
      __delay_data_791__delay_790__delay_789____variable_215 <= 0;
      __delay_data_792__delay_791__delay_790____variable_215 <= 0;
      __delay_data_793__delay_792__delay_791____variable_215 <= 0;
      _sra_data_233 <= 0;
      __variable_wdata_213 <= 0;
      __variable_wdata_214 <= 0;
      __variable_wdata_215 <= 0;
      _tmp_938 <= 0;
      _tmp_939 <= 0;
      _tmp_940 <= 0;
      _tmp_941 <= 0;
      _tmp_942 <= 0;
      _tmp_943 <= 0;
      _tmp_944 <= 0;
      _tmp_945 <= 0;
      _tmp_946 <= 0;
      _tmp_947 <= 0;
      _tmp_948 <= 0;
      _tmp_949 <= 0;
      _tmp_950 <= 0;
      _tmp_951 <= 0;
      _tmp_952 <= 0;
      _tmp_953 <= 0;
      _tmp_954 <= 0;
      _tmp_955 <= 0;
      _tmp_956 <= 0;
      _tmp_957 <= 0;
      _tmp_958 <= 0;
      _tmp_959 <= 0;
      _tmp_960 <= 0;
      _tmp_961 <= 0;
      _tmp_962 <= 0;
      _tmp_963 <= 0;
      _tmp_964 <= 0;
      _tmp_965 <= 0;
      _tmp_966 <= 0;
      _tmp_967 <= 0;
      _tmp_968 <= 0;
      _tmp_969 <= 0;
      _tmp_970 <= 0;
      _tmp_971 <= 0;
      _mul_10_busy_reg <= 0;
    end else begin
      if(_mul_10_stream_oready) begin
        _mul_10_x_source_ram_renable <= 0;
        _mul_10_x_source_fifo_deq <= 0;
      end 
      _mul_10_x_idle <= _mul_10_x_idle;
      if(_mul_10_stream_oready) begin
        _mul_10_y_source_ram_renable <= 0;
        _mul_10_y_source_fifo_deq <= 0;
      end 
      _mul_10_y_idle <= _mul_10_y_idle;
      if(_mul_10_stream_oready) begin
        _mul_10_rshift_source_ram_renable <= 0;
        _mul_10_rshift_source_fifo_deq <= 0;
      end 
      _mul_10_rshift_idle <= _mul_10_rshift_idle;
      if(_mul_10_stream_oready) begin
        _mul_10_z_sink_wenable <= 0;
        _mul_10_z_sink_fifo_enq <= 0;
      end 
      if(_mul_10_stream_oready) begin
        __mul_10_stream_ivalid_1 <= _mul_10_stream_ivalid;
      end 
      if(_mul_10_stream_oready) begin
        __mul_10_stream_ivalid_2 <= __mul_10_stream_ivalid_1;
      end 
      if(_mul_10_stream_oready) begin
        __mul_10_stream_ivalid_3 <= __mul_10_stream_ivalid_2;
      end 
      if(_mul_10_stream_oready) begin
        __mul_10_stream_ivalid_4 <= __mul_10_stream_ivalid_3;
      end 
      if(_mul_10_stream_oready) begin
        __mul_10_stream_ivalid_5 <= __mul_10_stream_ivalid_4;
      end 
      if(_mul_10_stream_oready) begin
        __mul_10_stream_ivalid_6 <= __mul_10_stream_ivalid_5;
      end 
      if(_mul_10_stream_oready) begin
        __mul_10_stream_ivalid_7 <= __mul_10_stream_ivalid_6;
      end 
      if(_mul_10_stream_oready) begin
        __mul_10_stream_ivalid_8 <= __mul_10_stream_ivalid_7;
      end 
      if(_mul_10_stream_oready) begin
        _greaterthan_data_216 <= mul_10_rshift_data > 1'sd0;
      end 
      if(_mul_10_stream_oready) begin
        _minus_data_218 <= mul_10_rshift_data - 2'sd1;
      end 
      if(_mul_10_stream_oready) begin
        _greatereq_data_229 <= mul_10_x_data >= 1'sd0;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_781__variable_213 <= mul_10_x_data;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_784__variable_214 <= mul_10_y_data;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_787__variable_215 <= mul_10_rshift_data;
      end 
      if(_mul_10_stream_oready) begin
        _sll_data_220 <= 2'sd1 << _minus_data_218;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_778_greaterthan_216 <= _greaterthan_data_216;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_779_greatereq_229 <= _greatereq_data_229;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_782__delay_781__variable_213 <= __delay_data_781__variable_213;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_785__delay_784__variable_214 <= __delay_data_784__variable_214;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_788__delay_787__variable_215 <= __delay_data_787__variable_215;
      end 
      if(_mul_10_stream_oready) begin
        _cond_data_226 <= (__delay_data_778_greaterthan_216)? _sll_data_220 : 1'sd0;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_780__delay_779_greatereq_229 <= __delay_data_779_greatereq_229;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_783__delay_782__delay_781__variable_213 <= __delay_data_782__delay_781__variable_213;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_786__delay_785__delay_784__variable_214 <= __delay_data_785__delay_784__variable_214;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_789__delay_788__delay_787__variable_215 <= __delay_data_788__delay_787__variable_215;
      end 
      if(_mul_10_stream_oready) begin
        __muladd_madd_odata_reg_232 <= __muladd_madd_odata_232;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_790__delay_789__delay_788____variable_215 <= __delay_data_789__delay_788__delay_787__variable_215;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_791__delay_790__delay_789____variable_215 <= __delay_data_790__delay_789__delay_788____variable_215;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_792__delay_791__delay_790____variable_215 <= __delay_data_791__delay_790__delay_789____variable_215;
      end 
      if(_mul_10_stream_oready) begin
        __delay_data_793__delay_792__delay_791____variable_215 <= __delay_data_792__delay_791__delay_790____variable_215;
      end 
      if(_mul_10_stream_oready) begin
        _sra_data_233 <= __muladd_data_232 >>> __delay_data_793__delay_792__delay_791____variable_215;
      end 
      if(__stream_conv2d_24_stream_ivalid_1 && _stream_conv2d_24_stream_oready) begin
        __variable_wdata_213 <= _cond_data_675;
      end 
      if(__stream_conv2d_24_stream_ivalid_1 && _stream_conv2d_24_stream_oready) begin
        __variable_wdata_214 <= __delay_data_1058_reinterpretcast_642;
      end 
      if(__stream_conv2d_24_stream_ivalid_1 && _stream_conv2d_24_stream_oready) begin
        __variable_wdata_215 <= _plus_data_794;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_938 <= _mul_10_source_start;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_939 <= _tmp_938;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_940 <= _tmp_939;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_941 <= _mul_10_source_start;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_942 <= _tmp_941;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_943 <= _tmp_942;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_944 <= _tmp_943;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_945 <= _tmp_944;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_946 <= _tmp_945;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_947 <= _tmp_946;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_948 <= _tmp_947;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_949 <= _tmp_948;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_950 <= _tmp_949;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_951 <= _mul_10_source_stop;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_952 <= _tmp_951;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_953 <= _tmp_952;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_954 <= _tmp_953;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_955 <= _tmp_954;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_956 <= _tmp_955;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_957 <= _tmp_956;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_958 <= _tmp_957;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_959 <= _tmp_958;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_960 <= _tmp_959;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_961 <= _mul_10_source_busy;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_962 <= _tmp_961;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_963 <= _tmp_962;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_964 <= _tmp_963;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_965 <= _tmp_964;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_966 <= _tmp_965;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_967 <= _tmp_966;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_968 <= _tmp_967;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_969 <= _tmp_968;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_970 <= _tmp_969;
      end 
      if(_mul_10_stream_oready) begin
        _tmp_971 <= _mul_10_sink_busy;
      end 
      if(!_mul_10_sink_busy && _tmp_971) begin
        _mul_10_busy_reg <= 0;
      end 
      if(_mul_10_source_busy) begin
        _mul_10_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_10_fsm_1 = 1;
  localparam _mul_10_fsm_2 = 2;
  localparam _mul_10_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_10_fsm <= _mul_10_fsm_init;
      _mul_10_source_start <= 0;
      _mul_10_source_busy <= 0;
      _mul_10_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_24_stream_ivalid_1 && _stream_conv2d_24_stream_oready) begin
        _mul_10_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_24_stream_oready && _stream_conv2d_24_busy) begin
        _mul_10_source_busy <= _stream_conv2d_24_source_busy;
      end 
      if(_mul_10_stream_oready && _tmp_940) begin
        _mul_10_stream_ivalid <= 1;
      end 
      if(_mul_10_stream_oready && 1'd0) begin
        _mul_10_stream_ivalid <= 0;
      end 
      case(_mul_10_fsm)
        _mul_10_fsm_init: begin
          if(_mul_10_run_flag) begin
            _mul_10_source_start <= 1;
          end 
          if(_mul_10_run_flag) begin
            _mul_10_fsm <= _mul_10_fsm_1;
          end 
        end
        _mul_10_fsm_1: begin
          if(_mul_10_source_start && _mul_10_stream_oready) begin
            _mul_10_source_start <= 0;
            _mul_10_source_busy <= 1;
          end 
          if(_mul_10_source_start && _mul_10_stream_oready) begin
            _mul_10_fsm <= _mul_10_fsm_2;
          end 
        end
        _mul_10_fsm_2: begin
          if(_mul_10_stream_oready) begin
            _mul_10_fsm <= _mul_10_fsm_3;
          end 
        end
        _mul_10_fsm_3: begin
          if(_mul_10_stream_oready && 1'd0) begin
            _mul_10_source_busy <= 0;
          end 
          if(_mul_10_stream_oready && 1'd0 && _mul_10_run_flag) begin
            _mul_10_source_start <= 1;
          end 
          if(_mul_10_stream_oready && 1'd0) begin
            _mul_10_fsm <= _mul_10_fsm_init;
          end 
          if(_mul_10_stream_oready && 1'd0 && _mul_10_run_flag) begin
            _mul_10_fsm <= _mul_10_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_11_x_source_ram_renable <= 0;
      _mul_11_x_source_fifo_deq <= 0;
      _mul_11_x_idle <= 1;
      _mul_11_y_source_ram_renable <= 0;
      _mul_11_y_source_fifo_deq <= 0;
      _mul_11_y_idle <= 1;
      _mul_11_rshift_source_ram_renable <= 0;
      _mul_11_rshift_source_fifo_deq <= 0;
      _mul_11_rshift_idle <= 1;
      _mul_11_z_sink_wenable <= 0;
      _mul_11_z_sink_fifo_enq <= 0;
      __mul_11_stream_ivalid_1 <= 0;
      __mul_11_stream_ivalid_2 <= 0;
      __mul_11_stream_ivalid_3 <= 0;
      __mul_11_stream_ivalid_4 <= 0;
      __mul_11_stream_ivalid_5 <= 0;
      __mul_11_stream_ivalid_6 <= 0;
      __mul_11_stream_ivalid_7 <= 0;
      __mul_11_stream_ivalid_8 <= 0;
      _greaterthan_data_237 <= 0;
      _minus_data_239 <= 0;
      _greatereq_data_250 <= 0;
      __delay_data_800__variable_234 <= 0;
      __delay_data_803__variable_235 <= 0;
      __delay_data_806__variable_236 <= 0;
      _sll_data_241 <= 0;
      __delay_data_797_greaterthan_237 <= 0;
      __delay_data_798_greatereq_250 <= 0;
      __delay_data_801__delay_800__variable_234 <= 0;
      __delay_data_804__delay_803__variable_235 <= 0;
      __delay_data_807__delay_806__variable_236 <= 0;
      _cond_data_247 <= 0;
      __delay_data_799__delay_798_greatereq_250 <= 0;
      __delay_data_802__delay_801__delay_800__variable_234 <= 0;
      __delay_data_805__delay_804__delay_803__variable_235 <= 0;
      __delay_data_808__delay_807__delay_806__variable_236 <= 0;
      __muladd_madd_odata_reg_253 <= 0;
      __delay_data_809__delay_808__delay_807____variable_236 <= 0;
      __delay_data_810__delay_809__delay_808____variable_236 <= 0;
      __delay_data_811__delay_810__delay_809____variable_236 <= 0;
      __delay_data_812__delay_811__delay_810____variable_236 <= 0;
      _sra_data_254 <= 0;
      __variable_wdata_234 <= 0;
      __variable_wdata_235 <= 0;
      __variable_wdata_236 <= 0;
      _tmp_972 <= 0;
      _tmp_973 <= 0;
      _tmp_974 <= 0;
      _tmp_975 <= 0;
      _tmp_976 <= 0;
      _tmp_977 <= 0;
      _tmp_978 <= 0;
      _tmp_979 <= 0;
      _tmp_980 <= 0;
      _tmp_981 <= 0;
      _tmp_982 <= 0;
      _tmp_983 <= 0;
      _tmp_984 <= 0;
      _tmp_985 <= 0;
      _tmp_986 <= 0;
      _tmp_987 <= 0;
      _tmp_988 <= 0;
      _tmp_989 <= 0;
      _tmp_990 <= 0;
      _tmp_991 <= 0;
      _tmp_992 <= 0;
      _tmp_993 <= 0;
      _tmp_994 <= 0;
      _tmp_995 <= 0;
      _tmp_996 <= 0;
      _tmp_997 <= 0;
      _tmp_998 <= 0;
      _tmp_999 <= 0;
      _tmp_1000 <= 0;
      _tmp_1001 <= 0;
      _tmp_1002 <= 0;
      _tmp_1003 <= 0;
      _tmp_1004 <= 0;
      _tmp_1005 <= 0;
      _mul_11_busy_reg <= 0;
    end else begin
      if(_mul_11_stream_oready) begin
        _mul_11_x_source_ram_renable <= 0;
        _mul_11_x_source_fifo_deq <= 0;
      end 
      _mul_11_x_idle <= _mul_11_x_idle;
      if(_mul_11_stream_oready) begin
        _mul_11_y_source_ram_renable <= 0;
        _mul_11_y_source_fifo_deq <= 0;
      end 
      _mul_11_y_idle <= _mul_11_y_idle;
      if(_mul_11_stream_oready) begin
        _mul_11_rshift_source_ram_renable <= 0;
        _mul_11_rshift_source_fifo_deq <= 0;
      end 
      _mul_11_rshift_idle <= _mul_11_rshift_idle;
      if(_mul_11_stream_oready) begin
        _mul_11_z_sink_wenable <= 0;
        _mul_11_z_sink_fifo_enq <= 0;
      end 
      if(_mul_11_stream_oready) begin
        __mul_11_stream_ivalid_1 <= _mul_11_stream_ivalid;
      end 
      if(_mul_11_stream_oready) begin
        __mul_11_stream_ivalid_2 <= __mul_11_stream_ivalid_1;
      end 
      if(_mul_11_stream_oready) begin
        __mul_11_stream_ivalid_3 <= __mul_11_stream_ivalid_2;
      end 
      if(_mul_11_stream_oready) begin
        __mul_11_stream_ivalid_4 <= __mul_11_stream_ivalid_3;
      end 
      if(_mul_11_stream_oready) begin
        __mul_11_stream_ivalid_5 <= __mul_11_stream_ivalid_4;
      end 
      if(_mul_11_stream_oready) begin
        __mul_11_stream_ivalid_6 <= __mul_11_stream_ivalid_5;
      end 
      if(_mul_11_stream_oready) begin
        __mul_11_stream_ivalid_7 <= __mul_11_stream_ivalid_6;
      end 
      if(_mul_11_stream_oready) begin
        __mul_11_stream_ivalid_8 <= __mul_11_stream_ivalid_7;
      end 
      if(_mul_11_stream_oready) begin
        _greaterthan_data_237 <= mul_11_rshift_data > 1'sd0;
      end 
      if(_mul_11_stream_oready) begin
        _minus_data_239 <= mul_11_rshift_data - 2'sd1;
      end 
      if(_mul_11_stream_oready) begin
        _greatereq_data_250 <= mul_11_x_data >= 1'sd0;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_800__variable_234 <= mul_11_x_data;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_803__variable_235 <= mul_11_y_data;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_806__variable_236 <= mul_11_rshift_data;
      end 
      if(_mul_11_stream_oready) begin
        _sll_data_241 <= 2'sd1 << _minus_data_239;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_797_greaterthan_237 <= _greaterthan_data_237;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_798_greatereq_250 <= _greatereq_data_250;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_801__delay_800__variable_234 <= __delay_data_800__variable_234;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_804__delay_803__variable_235 <= __delay_data_803__variable_235;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_807__delay_806__variable_236 <= __delay_data_806__variable_236;
      end 
      if(_mul_11_stream_oready) begin
        _cond_data_247 <= (__delay_data_797_greaterthan_237)? _sll_data_241 : 1'sd0;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_799__delay_798_greatereq_250 <= __delay_data_798_greatereq_250;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_802__delay_801__delay_800__variable_234 <= __delay_data_801__delay_800__variable_234;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_805__delay_804__delay_803__variable_235 <= __delay_data_804__delay_803__variable_235;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_808__delay_807__delay_806__variable_236 <= __delay_data_807__delay_806__variable_236;
      end 
      if(_mul_11_stream_oready) begin
        __muladd_madd_odata_reg_253 <= __muladd_madd_odata_253;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_809__delay_808__delay_807____variable_236 <= __delay_data_808__delay_807__delay_806__variable_236;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_810__delay_809__delay_808____variable_236 <= __delay_data_809__delay_808__delay_807____variable_236;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_811__delay_810__delay_809____variable_236 <= __delay_data_810__delay_809__delay_808____variable_236;
      end 
      if(_mul_11_stream_oready) begin
        __delay_data_812__delay_811__delay_810____variable_236 <= __delay_data_811__delay_810__delay_809____variable_236;
      end 
      if(_mul_11_stream_oready) begin
        _sra_data_254 <= __muladd_data_253 >>> __delay_data_812__delay_811__delay_810____variable_236;
      end 
      if(__stream_conv2d_24_stream_ivalid_1 && _stream_conv2d_24_stream_oready) begin
        __variable_wdata_234 <= _cond_data_677;
      end 
      if(__stream_conv2d_24_stream_ivalid_1 && _stream_conv2d_24_stream_oready) begin
        __variable_wdata_235 <= __delay_data_1060_reinterpretcast_643;
      end 
      if(__stream_conv2d_24_stream_ivalid_1 && _stream_conv2d_24_stream_oready) begin
        __variable_wdata_236 <= _plus_data_813;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_972 <= _mul_11_source_start;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_973 <= _tmp_972;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_974 <= _tmp_973;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_975 <= _mul_11_source_start;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_976 <= _tmp_975;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_977 <= _tmp_976;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_978 <= _tmp_977;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_979 <= _tmp_978;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_980 <= _tmp_979;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_981 <= _tmp_980;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_982 <= _tmp_981;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_983 <= _tmp_982;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_984 <= _tmp_983;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_985 <= _mul_11_source_stop;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_986 <= _tmp_985;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_987 <= _tmp_986;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_988 <= _tmp_987;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_989 <= _tmp_988;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_990 <= _tmp_989;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_991 <= _tmp_990;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_992 <= _tmp_991;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_993 <= _tmp_992;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_994 <= _tmp_993;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_995 <= _mul_11_source_busy;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_996 <= _tmp_995;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_997 <= _tmp_996;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_998 <= _tmp_997;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_999 <= _tmp_998;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_1000 <= _tmp_999;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_1001 <= _tmp_1000;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_1002 <= _tmp_1001;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_1003 <= _tmp_1002;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_1004 <= _tmp_1003;
      end 
      if(_mul_11_stream_oready) begin
        _tmp_1005 <= _mul_11_sink_busy;
      end 
      if(!_mul_11_sink_busy && _tmp_1005) begin
        _mul_11_busy_reg <= 0;
      end 
      if(_mul_11_source_busy) begin
        _mul_11_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_11_fsm_1 = 1;
  localparam _mul_11_fsm_2 = 2;
  localparam _mul_11_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_11_fsm <= _mul_11_fsm_init;
      _mul_11_source_start <= 0;
      _mul_11_source_busy <= 0;
      _mul_11_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_24_stream_ivalid_1 && _stream_conv2d_24_stream_oready) begin
        _mul_11_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_24_stream_oready && _stream_conv2d_24_busy) begin
        _mul_11_source_busy <= _stream_conv2d_24_source_busy;
      end 
      if(_mul_11_stream_oready && _tmp_974) begin
        _mul_11_stream_ivalid <= 1;
      end 
      if(_mul_11_stream_oready && 1'd0) begin
        _mul_11_stream_ivalid <= 0;
      end 
      case(_mul_11_fsm)
        _mul_11_fsm_init: begin
          if(_mul_11_run_flag) begin
            _mul_11_source_start <= 1;
          end 
          if(_mul_11_run_flag) begin
            _mul_11_fsm <= _mul_11_fsm_1;
          end 
        end
        _mul_11_fsm_1: begin
          if(_mul_11_source_start && _mul_11_stream_oready) begin
            _mul_11_source_start <= 0;
            _mul_11_source_busy <= 1;
          end 
          if(_mul_11_source_start && _mul_11_stream_oready) begin
            _mul_11_fsm <= _mul_11_fsm_2;
          end 
        end
        _mul_11_fsm_2: begin
          if(_mul_11_stream_oready) begin
            _mul_11_fsm <= _mul_11_fsm_3;
          end 
        end
        _mul_11_fsm_3: begin
          if(_mul_11_stream_oready && 1'd0) begin
            _mul_11_source_busy <= 0;
          end 
          if(_mul_11_stream_oready && 1'd0 && _mul_11_run_flag) begin
            _mul_11_source_start <= 1;
          end 
          if(_mul_11_stream_oready && 1'd0) begin
            _mul_11_fsm <= _mul_11_fsm_init;
          end 
          if(_mul_11_stream_oready && 1'd0 && _mul_11_run_flag) begin
            _mul_11_fsm <= _mul_11_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_12_x_source_ram_renable <= 0;
      _mul_12_x_source_fifo_deq <= 0;
      _mul_12_x_idle <= 1;
      _mul_12_y_source_ram_renable <= 0;
      _mul_12_y_source_fifo_deq <= 0;
      _mul_12_y_idle <= 1;
      _mul_12_rshift_source_ram_renable <= 0;
      _mul_12_rshift_source_fifo_deq <= 0;
      _mul_12_rshift_idle <= 1;
      _mul_12_z_sink_wenable <= 0;
      _mul_12_z_sink_fifo_enq <= 0;
      __mul_12_stream_ivalid_1 <= 0;
      __mul_12_stream_ivalid_2 <= 0;
      __mul_12_stream_ivalid_3 <= 0;
      __mul_12_stream_ivalid_4 <= 0;
      __mul_12_stream_ivalid_5 <= 0;
      __mul_12_stream_ivalid_6 <= 0;
      __mul_12_stream_ivalid_7 <= 0;
      __mul_12_stream_ivalid_8 <= 0;
      _greaterthan_data_258 <= 0;
      _minus_data_260 <= 0;
      _greatereq_data_271 <= 0;
      __delay_data_819__variable_255 <= 0;
      __delay_data_822__variable_256 <= 0;
      __delay_data_825__variable_257 <= 0;
      _sll_data_262 <= 0;
      __delay_data_816_greaterthan_258 <= 0;
      __delay_data_817_greatereq_271 <= 0;
      __delay_data_820__delay_819__variable_255 <= 0;
      __delay_data_823__delay_822__variable_256 <= 0;
      __delay_data_826__delay_825__variable_257 <= 0;
      _cond_data_268 <= 0;
      __delay_data_818__delay_817_greatereq_271 <= 0;
      __delay_data_821__delay_820__delay_819__variable_255 <= 0;
      __delay_data_824__delay_823__delay_822__variable_256 <= 0;
      __delay_data_827__delay_826__delay_825__variable_257 <= 0;
      __muladd_madd_odata_reg_274 <= 0;
      __delay_data_828__delay_827__delay_826____variable_257 <= 0;
      __delay_data_829__delay_828__delay_827____variable_257 <= 0;
      __delay_data_830__delay_829__delay_828____variable_257 <= 0;
      __delay_data_831__delay_830__delay_829____variable_257 <= 0;
      _sra_data_275 <= 0;
      __variable_wdata_255 <= 0;
      __variable_wdata_256 <= 0;
      __variable_wdata_257 <= 0;
      _tmp_1006 <= 0;
      _tmp_1007 <= 0;
      _tmp_1008 <= 0;
      _tmp_1009 <= 0;
      _tmp_1010 <= 0;
      _tmp_1011 <= 0;
      _tmp_1012 <= 0;
      _tmp_1013 <= 0;
      _tmp_1014 <= 0;
      _tmp_1015 <= 0;
      _tmp_1016 <= 0;
      _tmp_1017 <= 0;
      _tmp_1018 <= 0;
      _tmp_1019 <= 0;
      _tmp_1020 <= 0;
      _tmp_1021 <= 0;
      _tmp_1022 <= 0;
      _tmp_1023 <= 0;
      _tmp_1024 <= 0;
      _tmp_1025 <= 0;
      _tmp_1026 <= 0;
      _tmp_1027 <= 0;
      _tmp_1028 <= 0;
      _tmp_1029 <= 0;
      _tmp_1030 <= 0;
      _tmp_1031 <= 0;
      _tmp_1032 <= 0;
      _tmp_1033 <= 0;
      _tmp_1034 <= 0;
      _tmp_1035 <= 0;
      _tmp_1036 <= 0;
      _tmp_1037 <= 0;
      _tmp_1038 <= 0;
      _tmp_1039 <= 0;
      _mul_12_busy_reg <= 0;
    end else begin
      if(_mul_12_stream_oready) begin
        _mul_12_x_source_ram_renable <= 0;
        _mul_12_x_source_fifo_deq <= 0;
      end 
      _mul_12_x_idle <= _mul_12_x_idle;
      if(_mul_12_stream_oready) begin
        _mul_12_y_source_ram_renable <= 0;
        _mul_12_y_source_fifo_deq <= 0;
      end 
      _mul_12_y_idle <= _mul_12_y_idle;
      if(_mul_12_stream_oready) begin
        _mul_12_rshift_source_ram_renable <= 0;
        _mul_12_rshift_source_fifo_deq <= 0;
      end 
      _mul_12_rshift_idle <= _mul_12_rshift_idle;
      if(_mul_12_stream_oready) begin
        _mul_12_z_sink_wenable <= 0;
        _mul_12_z_sink_fifo_enq <= 0;
      end 
      if(_mul_12_stream_oready) begin
        __mul_12_stream_ivalid_1 <= _mul_12_stream_ivalid;
      end 
      if(_mul_12_stream_oready) begin
        __mul_12_stream_ivalid_2 <= __mul_12_stream_ivalid_1;
      end 
      if(_mul_12_stream_oready) begin
        __mul_12_stream_ivalid_3 <= __mul_12_stream_ivalid_2;
      end 
      if(_mul_12_stream_oready) begin
        __mul_12_stream_ivalid_4 <= __mul_12_stream_ivalid_3;
      end 
      if(_mul_12_stream_oready) begin
        __mul_12_stream_ivalid_5 <= __mul_12_stream_ivalid_4;
      end 
      if(_mul_12_stream_oready) begin
        __mul_12_stream_ivalid_6 <= __mul_12_stream_ivalid_5;
      end 
      if(_mul_12_stream_oready) begin
        __mul_12_stream_ivalid_7 <= __mul_12_stream_ivalid_6;
      end 
      if(_mul_12_stream_oready) begin
        __mul_12_stream_ivalid_8 <= __mul_12_stream_ivalid_7;
      end 
      if(_mul_12_stream_oready) begin
        _greaterthan_data_258 <= mul_12_rshift_data > 1'sd0;
      end 
      if(_mul_12_stream_oready) begin
        _minus_data_260 <= mul_12_rshift_data - 2'sd1;
      end 
      if(_mul_12_stream_oready) begin
        _greatereq_data_271 <= mul_12_x_data >= 1'sd0;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_819__variable_255 <= mul_12_x_data;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_822__variable_256 <= mul_12_y_data;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_825__variable_257 <= mul_12_rshift_data;
      end 
      if(_mul_12_stream_oready) begin
        _sll_data_262 <= 2'sd1 << _minus_data_260;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_816_greaterthan_258 <= _greaterthan_data_258;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_817_greatereq_271 <= _greatereq_data_271;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_820__delay_819__variable_255 <= __delay_data_819__variable_255;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_823__delay_822__variable_256 <= __delay_data_822__variable_256;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_826__delay_825__variable_257 <= __delay_data_825__variable_257;
      end 
      if(_mul_12_stream_oready) begin
        _cond_data_268 <= (__delay_data_816_greaterthan_258)? _sll_data_262 : 1'sd0;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_818__delay_817_greatereq_271 <= __delay_data_817_greatereq_271;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_821__delay_820__delay_819__variable_255 <= __delay_data_820__delay_819__variable_255;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_824__delay_823__delay_822__variable_256 <= __delay_data_823__delay_822__variable_256;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_827__delay_826__delay_825__variable_257 <= __delay_data_826__delay_825__variable_257;
      end 
      if(_mul_12_stream_oready) begin
        __muladd_madd_odata_reg_274 <= __muladd_madd_odata_274;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_828__delay_827__delay_826____variable_257 <= __delay_data_827__delay_826__delay_825__variable_257;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_829__delay_828__delay_827____variable_257 <= __delay_data_828__delay_827__delay_826____variable_257;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_830__delay_829__delay_828____variable_257 <= __delay_data_829__delay_828__delay_827____variable_257;
      end 
      if(_mul_12_stream_oready) begin
        __delay_data_831__delay_830__delay_829____variable_257 <= __delay_data_830__delay_829__delay_828____variable_257;
      end 
      if(_mul_12_stream_oready) begin
        _sra_data_275 <= __muladd_data_274 >>> __delay_data_831__delay_830__delay_829____variable_257;
      end 
      if(__stream_conv2d_24_stream_ivalid_1 && _stream_conv2d_24_stream_oready) begin
        __variable_wdata_255 <= _cond_data_679;
      end 
      if(__stream_conv2d_24_stream_ivalid_1 && _stream_conv2d_24_stream_oready) begin
        __variable_wdata_256 <= __delay_data_1062_reinterpretcast_644;
      end 
      if(__stream_conv2d_24_stream_ivalid_1 && _stream_conv2d_24_stream_oready) begin
        __variable_wdata_257 <= _plus_data_832;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_1006 <= _mul_12_source_start;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_1007 <= _tmp_1006;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_1008 <= _tmp_1007;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_1009 <= _mul_12_source_start;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_1010 <= _tmp_1009;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_1011 <= _tmp_1010;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_1012 <= _tmp_1011;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_1013 <= _tmp_1012;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_1014 <= _tmp_1013;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_1015 <= _tmp_1014;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_1016 <= _tmp_1015;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_1017 <= _tmp_1016;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_1018 <= _tmp_1017;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_1019 <= _mul_12_source_stop;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_1020 <= _tmp_1019;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_1021 <= _tmp_1020;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_1022 <= _tmp_1021;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_1023 <= _tmp_1022;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_1024 <= _tmp_1023;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_1025 <= _tmp_1024;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_1026 <= _tmp_1025;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_1027 <= _tmp_1026;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_1028 <= _tmp_1027;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_1029 <= _mul_12_source_busy;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_1030 <= _tmp_1029;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_1031 <= _tmp_1030;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_1032 <= _tmp_1031;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_1033 <= _tmp_1032;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_1034 <= _tmp_1033;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_1035 <= _tmp_1034;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_1036 <= _tmp_1035;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_1037 <= _tmp_1036;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_1038 <= _tmp_1037;
      end 
      if(_mul_12_stream_oready) begin
        _tmp_1039 <= _mul_12_sink_busy;
      end 
      if(!_mul_12_sink_busy && _tmp_1039) begin
        _mul_12_busy_reg <= 0;
      end 
      if(_mul_12_source_busy) begin
        _mul_12_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_12_fsm_1 = 1;
  localparam _mul_12_fsm_2 = 2;
  localparam _mul_12_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_12_fsm <= _mul_12_fsm_init;
      _mul_12_source_start <= 0;
      _mul_12_source_busy <= 0;
      _mul_12_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_24_stream_ivalid_1 && _stream_conv2d_24_stream_oready) begin
        _mul_12_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_24_stream_oready && _stream_conv2d_24_busy) begin
        _mul_12_source_busy <= _stream_conv2d_24_source_busy;
      end 
      if(_mul_12_stream_oready && _tmp_1008) begin
        _mul_12_stream_ivalid <= 1;
      end 
      if(_mul_12_stream_oready && 1'd0) begin
        _mul_12_stream_ivalid <= 0;
      end 
      case(_mul_12_fsm)
        _mul_12_fsm_init: begin
          if(_mul_12_run_flag) begin
            _mul_12_source_start <= 1;
          end 
          if(_mul_12_run_flag) begin
            _mul_12_fsm <= _mul_12_fsm_1;
          end 
        end
        _mul_12_fsm_1: begin
          if(_mul_12_source_start && _mul_12_stream_oready) begin
            _mul_12_source_start <= 0;
            _mul_12_source_busy <= 1;
          end 
          if(_mul_12_source_start && _mul_12_stream_oready) begin
            _mul_12_fsm <= _mul_12_fsm_2;
          end 
        end
        _mul_12_fsm_2: begin
          if(_mul_12_stream_oready) begin
            _mul_12_fsm <= _mul_12_fsm_3;
          end 
        end
        _mul_12_fsm_3: begin
          if(_mul_12_stream_oready && 1'd0) begin
            _mul_12_source_busy <= 0;
          end 
          if(_mul_12_stream_oready && 1'd0 && _mul_12_run_flag) begin
            _mul_12_source_start <= 1;
          end 
          if(_mul_12_stream_oready && 1'd0) begin
            _mul_12_fsm <= _mul_12_fsm_init;
          end 
          if(_mul_12_stream_oready && 1'd0 && _mul_12_run_flag) begin
            _mul_12_fsm <= _mul_12_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_13_x_source_ram_renable <= 0;
      _mul_13_x_source_fifo_deq <= 0;
      _mul_13_x_idle <= 1;
      _mul_13_y_source_ram_renable <= 0;
      _mul_13_y_source_fifo_deq <= 0;
      _mul_13_y_idle <= 1;
      _mul_13_rshift_source_ram_renable <= 0;
      _mul_13_rshift_source_fifo_deq <= 0;
      _mul_13_rshift_idle <= 1;
      _mul_13_z_sink_wenable <= 0;
      _mul_13_z_sink_fifo_enq <= 0;
      __mul_13_stream_ivalid_1 <= 0;
      __mul_13_stream_ivalid_2 <= 0;
      __mul_13_stream_ivalid_3 <= 0;
      __mul_13_stream_ivalid_4 <= 0;
      __mul_13_stream_ivalid_5 <= 0;
      __mul_13_stream_ivalid_6 <= 0;
      __mul_13_stream_ivalid_7 <= 0;
      __mul_13_stream_ivalid_8 <= 0;
      _greaterthan_data_279 <= 0;
      _minus_data_281 <= 0;
      _greatereq_data_292 <= 0;
      __delay_data_838__variable_276 <= 0;
      __delay_data_841__variable_277 <= 0;
      __delay_data_844__variable_278 <= 0;
      _sll_data_283 <= 0;
      __delay_data_835_greaterthan_279 <= 0;
      __delay_data_836_greatereq_292 <= 0;
      __delay_data_839__delay_838__variable_276 <= 0;
      __delay_data_842__delay_841__variable_277 <= 0;
      __delay_data_845__delay_844__variable_278 <= 0;
      _cond_data_289 <= 0;
      __delay_data_837__delay_836_greatereq_292 <= 0;
      __delay_data_840__delay_839__delay_838__variable_276 <= 0;
      __delay_data_843__delay_842__delay_841__variable_277 <= 0;
      __delay_data_846__delay_845__delay_844__variable_278 <= 0;
      __muladd_madd_odata_reg_295 <= 0;
      __delay_data_847__delay_846__delay_845____variable_278 <= 0;
      __delay_data_848__delay_847__delay_846____variable_278 <= 0;
      __delay_data_849__delay_848__delay_847____variable_278 <= 0;
      __delay_data_850__delay_849__delay_848____variable_278 <= 0;
      _sra_data_296 <= 0;
      __variable_wdata_276 <= 0;
      __variable_wdata_277 <= 0;
      __variable_wdata_278 <= 0;
      _tmp_1040 <= 0;
      _tmp_1041 <= 0;
      _tmp_1042 <= 0;
      _tmp_1043 <= 0;
      _tmp_1044 <= 0;
      _tmp_1045 <= 0;
      _tmp_1046 <= 0;
      _tmp_1047 <= 0;
      _tmp_1048 <= 0;
      _tmp_1049 <= 0;
      _tmp_1050 <= 0;
      _tmp_1051 <= 0;
      _tmp_1052 <= 0;
      _tmp_1053 <= 0;
      _tmp_1054 <= 0;
      _tmp_1055 <= 0;
      _tmp_1056 <= 0;
      _tmp_1057 <= 0;
      _tmp_1058 <= 0;
      _tmp_1059 <= 0;
      _tmp_1060 <= 0;
      _tmp_1061 <= 0;
      _tmp_1062 <= 0;
      _tmp_1063 <= 0;
      _tmp_1064 <= 0;
      _tmp_1065 <= 0;
      _tmp_1066 <= 0;
      _tmp_1067 <= 0;
      _tmp_1068 <= 0;
      _tmp_1069 <= 0;
      _tmp_1070 <= 0;
      _tmp_1071 <= 0;
      _tmp_1072 <= 0;
      _tmp_1073 <= 0;
      _mul_13_busy_reg <= 0;
    end else begin
      if(_mul_13_stream_oready) begin
        _mul_13_x_source_ram_renable <= 0;
        _mul_13_x_source_fifo_deq <= 0;
      end 
      _mul_13_x_idle <= _mul_13_x_idle;
      if(_mul_13_stream_oready) begin
        _mul_13_y_source_ram_renable <= 0;
        _mul_13_y_source_fifo_deq <= 0;
      end 
      _mul_13_y_idle <= _mul_13_y_idle;
      if(_mul_13_stream_oready) begin
        _mul_13_rshift_source_ram_renable <= 0;
        _mul_13_rshift_source_fifo_deq <= 0;
      end 
      _mul_13_rshift_idle <= _mul_13_rshift_idle;
      if(_mul_13_stream_oready) begin
        _mul_13_z_sink_wenable <= 0;
        _mul_13_z_sink_fifo_enq <= 0;
      end 
      if(_mul_13_stream_oready) begin
        __mul_13_stream_ivalid_1 <= _mul_13_stream_ivalid;
      end 
      if(_mul_13_stream_oready) begin
        __mul_13_stream_ivalid_2 <= __mul_13_stream_ivalid_1;
      end 
      if(_mul_13_stream_oready) begin
        __mul_13_stream_ivalid_3 <= __mul_13_stream_ivalid_2;
      end 
      if(_mul_13_stream_oready) begin
        __mul_13_stream_ivalid_4 <= __mul_13_stream_ivalid_3;
      end 
      if(_mul_13_stream_oready) begin
        __mul_13_stream_ivalid_5 <= __mul_13_stream_ivalid_4;
      end 
      if(_mul_13_stream_oready) begin
        __mul_13_stream_ivalid_6 <= __mul_13_stream_ivalid_5;
      end 
      if(_mul_13_stream_oready) begin
        __mul_13_stream_ivalid_7 <= __mul_13_stream_ivalid_6;
      end 
      if(_mul_13_stream_oready) begin
        __mul_13_stream_ivalid_8 <= __mul_13_stream_ivalid_7;
      end 
      if(_mul_13_stream_oready) begin
        _greaterthan_data_279 <= mul_13_rshift_data > 1'sd0;
      end 
      if(_mul_13_stream_oready) begin
        _minus_data_281 <= mul_13_rshift_data - 2'sd1;
      end 
      if(_mul_13_stream_oready) begin
        _greatereq_data_292 <= mul_13_x_data >= 1'sd0;
      end 
      if(_mul_13_stream_oready) begin
        __delay_data_838__variable_276 <= mul_13_x_data;
      end 
      if(_mul_13_stream_oready) begin
        __delay_data_841__variable_277 <= mul_13_y_data;
      end 
      if(_mul_13_stream_oready) begin
        __delay_data_844__variable_278 <= mul_13_rshift_data;
      end 
      if(_mul_13_stream_oready) begin
        _sll_data_283 <= 2'sd1 << _minus_data_281;
      end 
      if(_mul_13_stream_oready) begin
        __delay_data_835_greaterthan_279 <= _greaterthan_data_279;
      end 
      if(_mul_13_stream_oready) begin
        __delay_data_836_greatereq_292 <= _greatereq_data_292;
      end 
      if(_mul_13_stream_oready) begin
        __delay_data_839__delay_838__variable_276 <= __delay_data_838__variable_276;
      end 
      if(_mul_13_stream_oready) begin
        __delay_data_842__delay_841__variable_277 <= __delay_data_841__variable_277;
      end 
      if(_mul_13_stream_oready) begin
        __delay_data_845__delay_844__variable_278 <= __delay_data_844__variable_278;
      end 
      if(_mul_13_stream_oready) begin
        _cond_data_289 <= (__delay_data_835_greaterthan_279)? _sll_data_283 : 1'sd0;
      end 
      if(_mul_13_stream_oready) begin
        __delay_data_837__delay_836_greatereq_292 <= __delay_data_836_greatereq_292;
      end 
      if(_mul_13_stream_oready) begin
        __delay_data_840__delay_839__delay_838__variable_276 <= __delay_data_839__delay_838__variable_276;
      end 
      if(_mul_13_stream_oready) begin
        __delay_data_843__delay_842__delay_841__variable_277 <= __delay_data_842__delay_841__variable_277;
      end 
      if(_mul_13_stream_oready) begin
        __delay_data_846__delay_845__delay_844__variable_278 <= __delay_data_845__delay_844__variable_278;
      end 
      if(_mul_13_stream_oready) begin
        __muladd_madd_odata_reg_295 <= __muladd_madd_odata_295;
      end 
      if(_mul_13_stream_oready) begin
        __delay_data_847__delay_846__delay_845____variable_278 <= __delay_data_846__delay_845__delay_844__variable_278;
      end 
      if(_mul_13_stream_oready) begin
        __delay_data_848__delay_847__delay_846____variable_278 <= __delay_data_847__delay_846__delay_845____variable_278;
      end 
      if(_mul_13_stream_oready) begin
        __delay_data_849__delay_848__delay_847____variable_278 <= __delay_data_848__delay_847__delay_846____variable_278;
      end 
      if(_mul_13_stream_oready) begin
        __delay_data_850__delay_849__delay_848____variable_278 <= __delay_data_849__delay_848__delay_847____variable_278;
      end 
      if(_mul_13_stream_oready) begin
        _sra_data_296 <= __muladd_data_295 >>> __delay_data_850__delay_849__delay_848____variable_278;
      end 
      if(__stream_conv2d_24_stream_ivalid_1 && _stream_conv2d_24_stream_oready) begin
        __variable_wdata_276 <= _cond_data_681;
      end 
      if(__stream_conv2d_24_stream_ivalid_1 && _stream_conv2d_24_stream_oready) begin
        __variable_wdata_277 <= __delay_data_1064_reinterpretcast_645;
      end 
      if(__stream_conv2d_24_stream_ivalid_1 && _stream_conv2d_24_stream_oready) begin
        __variable_wdata_278 <= _plus_data_851;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_1040 <= _mul_13_source_start;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_1041 <= _tmp_1040;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_1042 <= _tmp_1041;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_1043 <= _mul_13_source_start;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_1044 <= _tmp_1043;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_1045 <= _tmp_1044;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_1046 <= _tmp_1045;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_1047 <= _tmp_1046;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_1048 <= _tmp_1047;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_1049 <= _tmp_1048;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_1050 <= _tmp_1049;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_1051 <= _tmp_1050;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_1052 <= _tmp_1051;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_1053 <= _mul_13_source_stop;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_1054 <= _tmp_1053;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_1055 <= _tmp_1054;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_1056 <= _tmp_1055;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_1057 <= _tmp_1056;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_1058 <= _tmp_1057;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_1059 <= _tmp_1058;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_1060 <= _tmp_1059;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_1061 <= _tmp_1060;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_1062 <= _tmp_1061;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_1063 <= _mul_13_source_busy;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_1064 <= _tmp_1063;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_1065 <= _tmp_1064;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_1066 <= _tmp_1065;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_1067 <= _tmp_1066;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_1068 <= _tmp_1067;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_1069 <= _tmp_1068;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_1070 <= _tmp_1069;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_1071 <= _tmp_1070;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_1072 <= _tmp_1071;
      end 
      if(_mul_13_stream_oready) begin
        _tmp_1073 <= _mul_13_sink_busy;
      end 
      if(!_mul_13_sink_busy && _tmp_1073) begin
        _mul_13_busy_reg <= 0;
      end 
      if(_mul_13_source_busy) begin
        _mul_13_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_13_fsm_1 = 1;
  localparam _mul_13_fsm_2 = 2;
  localparam _mul_13_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_13_fsm <= _mul_13_fsm_init;
      _mul_13_source_start <= 0;
      _mul_13_source_busy <= 0;
      _mul_13_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_24_stream_ivalid_1 && _stream_conv2d_24_stream_oready) begin
        _mul_13_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_24_stream_oready && _stream_conv2d_24_busy) begin
        _mul_13_source_busy <= _stream_conv2d_24_source_busy;
      end 
      if(_mul_13_stream_oready && _tmp_1042) begin
        _mul_13_stream_ivalid <= 1;
      end 
      if(_mul_13_stream_oready && 1'd0) begin
        _mul_13_stream_ivalid <= 0;
      end 
      case(_mul_13_fsm)
        _mul_13_fsm_init: begin
          if(_mul_13_run_flag) begin
            _mul_13_source_start <= 1;
          end 
          if(_mul_13_run_flag) begin
            _mul_13_fsm <= _mul_13_fsm_1;
          end 
        end
        _mul_13_fsm_1: begin
          if(_mul_13_source_start && _mul_13_stream_oready) begin
            _mul_13_source_start <= 0;
            _mul_13_source_busy <= 1;
          end 
          if(_mul_13_source_start && _mul_13_stream_oready) begin
            _mul_13_fsm <= _mul_13_fsm_2;
          end 
        end
        _mul_13_fsm_2: begin
          if(_mul_13_stream_oready) begin
            _mul_13_fsm <= _mul_13_fsm_3;
          end 
        end
        _mul_13_fsm_3: begin
          if(_mul_13_stream_oready && 1'd0) begin
            _mul_13_source_busy <= 0;
          end 
          if(_mul_13_stream_oready && 1'd0 && _mul_13_run_flag) begin
            _mul_13_source_start <= 1;
          end 
          if(_mul_13_stream_oready && 1'd0) begin
            _mul_13_fsm <= _mul_13_fsm_init;
          end 
          if(_mul_13_stream_oready && 1'd0 && _mul_13_run_flag) begin
            _mul_13_fsm <= _mul_13_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __reduce_max_14_x_source_ram_renable <= 0;
      __reduce_max_14_x_source_fifo_deq <= 0;
      __reduce_max_14_x_idle <= 1;
      __reduce_max_14_data_sink_wenable <= 0;
      __reduce_max_14_data_sink_fifo_enq <= 0;
      __reduce_max_14_valid_sink_wenable <= 0;
      __reduce_max_14_valid_sink_fifo_enq <= 0;
      ___reduce_max_14_stream_ivalid_1 <= 0;
      _reducemax_data_300 <= -9'sd128;
      _reducemax_count_300 <= 0;
      _reducemax_prev_count_max_300 <= 0;
      _pulse_data_302 <= 1'sd0;
      _pulse_count_302 <= 0;
      _pulse_prev_count_max_302 <= 0;
      __variable_wdata_299 <= 0;
      __variable_wdata_297 <= 0;
      __variable_wdata_298 <= 0;
      _tmp_1390 <= 0;
      _tmp_1391 <= 0;
      _tmp_1392 <= 0;
      _tmp_1393 <= 0;
      _tmp_1394 <= 0;
      _tmp_1395 <= 0;
      _tmp_1396 <= 0;
      _tmp_1397 <= 0;
      _tmp_1398 <= 0;
      _tmp_1399 <= 0;
      _tmp_1400 <= 0;
      _tmp_1401 <= 0;
      _tmp_1402 <= 0;
      _tmp_1403 <= 0;
      _tmp_1404 <= 0;
      _tmp_1405 <= 0;
      _tmp_1406 <= 0;
      _tmp_1407 <= 0;
      _tmp_1408 <= 0;
      _tmp_1409 <= 0;
      __reduce_max_14_busy_reg <= 0;
    end else begin
      if(__reduce_max_14_stream_oready) begin
        __reduce_max_14_x_source_ram_renable <= 0;
        __reduce_max_14_x_source_fifo_deq <= 0;
      end 
      __reduce_max_14_x_idle <= __reduce_max_14_x_idle;
      if(__reduce_max_14_stream_oready) begin
        __reduce_max_14_data_sink_wenable <= 0;
        __reduce_max_14_data_sink_fifo_enq <= 0;
      end 
      if(__reduce_max_14_stream_oready) begin
        __reduce_max_14_valid_sink_wenable <= 0;
        __reduce_max_14_valid_sink_fifo_enq <= 0;
      end 
      if(__reduce_max_14_stream_oready) begin
        ___reduce_max_14_stream_ivalid_1 <= __reduce_max_14_stream_ivalid;
      end 
      if(__reduce_max_14_stream_ivalid && __reduce_max_14_stream_oready && _reducemax_reset_cond_300) begin
        _reducemax_data_300 <= -9'sd128;
      end 
      if(__reduce_max_14_stream_ivalid && __reduce_max_14_stream_oready) begin
        _reducemax_count_300 <= (_reducemax_current_count_300 >= _reduce_max_14_size_data - 1)? 0 : _reducemax_current_count_300 + 1;
      end 
      if(__reduce_max_14_stream_ivalid && __reduce_max_14_stream_oready) begin
        _reducemax_prev_count_max_300 <= _reducemax_current_count_300 >= _reduce_max_14_size_data - 1;
      end 
      if(__reduce_max_14_stream_ivalid && __reduce_max_14_stream_oready) begin
        _reducemax_data_300 <= (_reducemax_current_data_300 < _reduce_max_14_x_data)? _reduce_max_14_x_data : _reducemax_current_data_300;
      end 
      if(__reduce_max_14_stream_ivalid && __reduce_max_14_stream_oready && _pulse_reset_cond_302) begin
        _pulse_data_302 <= 1'sd0;
      end 
      if(__reduce_max_14_stream_ivalid && __reduce_max_14_stream_oready) begin
        _pulse_count_302 <= (_pulse_current_count_302 >= _reduce_max_14_size_data - 1)? 0 : _pulse_current_count_302 + 1;
      end 
      if(__reduce_max_14_stream_ivalid && __reduce_max_14_stream_oready) begin
        _pulse_prev_count_max_302 <= _pulse_current_count_302 >= _reduce_max_14_size_data - 1;
      end 
      if(__reduce_max_14_stream_ivalid && __reduce_max_14_stream_oready) begin
        _pulse_data_302 <= _pulse_current_count_302 >= _reduce_max_14_size_data - 1;
      end 
      if(__stream_max_pool_serial_26_stream_ivalid_3 && _stream_max_pool_serial_26_stream_oready) begin
        __variable_wdata_299 <= __delay_data_1179__delay_1178__delay_1177__variable_896;
      end 
      if(__stream_max_pool_serial_26_stream_ivalid_3 && _stream_max_pool_serial_26_stream_oready) begin
        __variable_wdata_297 <= _cond_data_907;
      end 
      if(__stream_max_pool_serial_26_stream_ivalid_3 && _stream_max_pool_serial_26_stream_oready) begin
        __variable_wdata_298 <= __delay_data_1182__delay_1181__delay_1180__variable_893;
      end 
      if(__reduce_max_14_stream_oready) begin
        _tmp_1390 <= __reduce_max_14_source_start;
      end 
      if(__reduce_max_14_stream_oready) begin
        _tmp_1391 <= _tmp_1390;
      end 
      if(__reduce_max_14_stream_oready) begin
        _tmp_1392 <= _tmp_1391;
      end 
      if(__reduce_max_14_stream_oready) begin
        _tmp_1393 <= __reduce_max_14_source_start;
      end 
      if(__reduce_max_14_stream_oready) begin
        _tmp_1394 <= _tmp_1393;
      end 
      if(__reduce_max_14_stream_oready) begin
        _tmp_1395 <= _tmp_1394;
      end 
      if(__reduce_max_14_stream_oready && _tmp_1395) begin
        __variable_wdata_299 <= 1;
      end 
      if(__reduce_max_14_stream_oready) begin
        _tmp_1396 <= __reduce_max_14_source_start;
      end 
      if(__reduce_max_14_stream_oready) begin
        _tmp_1397 <= _tmp_1396;
      end 
      if(__reduce_max_14_stream_oready) begin
        _tmp_1398 <= _tmp_1397;
      end 
      if(__reduce_max_14_stream_oready) begin
        _tmp_1399 <= _tmp_1398;
      end 
      if(__reduce_max_14_stream_oready && _tmp_1399) begin
        __variable_wdata_299 <= 0;
      end 
      if(__reduce_max_14_stream_oready && 1'd0) begin
        __variable_wdata_299 <= 1;
      end 
      if(__reduce_max_14_stream_oready) begin
        _tmp_1400 <= __reduce_max_14_source_start;
      end 
      if(__reduce_max_14_stream_oready) begin
        _tmp_1401 <= _tmp_1400;
      end 
      if(__reduce_max_14_stream_oready) begin
        _tmp_1402 <= _tmp_1401;
      end 
      if(__reduce_max_14_stream_oready) begin
        _tmp_1403 <= __reduce_max_14_source_stop;
      end 
      if(__reduce_max_14_stream_oready) begin
        _tmp_1404 <= _tmp_1403;
      end 
      if(__reduce_max_14_stream_oready) begin
        _tmp_1405 <= _tmp_1404;
      end 
      if(__reduce_max_14_stream_oready) begin
        _tmp_1406 <= __reduce_max_14_source_busy;
      end 
      if(__reduce_max_14_stream_oready) begin
        _tmp_1407 <= _tmp_1406;
      end 
      if(__reduce_max_14_stream_oready) begin
        _tmp_1408 <= _tmp_1407;
      end 
      if(__reduce_max_14_stream_oready) begin
        _tmp_1409 <= __reduce_max_14_sink_busy;
      end 
      if(!__reduce_max_14_sink_busy && _tmp_1409) begin
        __reduce_max_14_busy_reg <= 0;
      end 
      if(__reduce_max_14_source_busy) begin
        __reduce_max_14_busy_reg <= 1;
      end 
    end
  end

  localparam __reduce_max_14_fsm_1 = 1;
  localparam __reduce_max_14_fsm_2 = 2;
  localparam __reduce_max_14_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      __reduce_max_14_fsm <= __reduce_max_14_fsm_init;
      __reduce_max_14_source_start <= 0;
      __reduce_max_14_source_busy <= 0;
      __reduce_max_14_stream_ivalid <= 0;
    end else begin
      if(__stream_max_pool_serial_26_stream_ivalid_3 && _stream_max_pool_serial_26_stream_oready) begin
        __reduce_max_14_stream_ivalid <= 1'd1;
      end 
      if(_stream_max_pool_serial_26_stream_oready && _stream_max_pool_serial_26_busy) begin
        __reduce_max_14_source_busy <= _stream_max_pool_serial_26_source_busy;
      end 
      if(__reduce_max_14_stream_oready && _tmp_1392) begin
        __reduce_max_14_stream_ivalid <= 1;
      end 
      if(__reduce_max_14_stream_oready && 1'd0) begin
        __reduce_max_14_stream_ivalid <= 0;
      end 
      case(__reduce_max_14_fsm)
        __reduce_max_14_fsm_init: begin
          if(__reduce_max_14_run_flag) begin
            __reduce_max_14_source_start <= 1;
          end 
          if(__reduce_max_14_run_flag) begin
            __reduce_max_14_fsm <= __reduce_max_14_fsm_1;
          end 
        end
        __reduce_max_14_fsm_1: begin
          if(__reduce_max_14_source_start && __reduce_max_14_stream_oready) begin
            __reduce_max_14_source_start <= 0;
            __reduce_max_14_source_busy <= 1;
          end 
          if(__reduce_max_14_source_start && __reduce_max_14_stream_oready) begin
            __reduce_max_14_fsm <= __reduce_max_14_fsm_2;
          end 
        end
        __reduce_max_14_fsm_2: begin
          if(__reduce_max_14_stream_oready) begin
            __reduce_max_14_fsm <= __reduce_max_14_fsm_3;
          end 
        end
        __reduce_max_14_fsm_3: begin
          if(__reduce_max_14_stream_oready && 1'd0) begin
            __reduce_max_14_source_busy <= 0;
          end 
          if(__reduce_max_14_stream_oready && 1'd0 && __reduce_max_14_run_flag) begin
            __reduce_max_14_source_start <= 1;
          end 
          if(__reduce_max_14_stream_oready && 1'd0) begin
            __reduce_max_14_fsm <= __reduce_max_14_fsm_init;
          end 
          if(__reduce_max_14_stream_oready && 1'd0 && __reduce_max_14_run_flag) begin
            __reduce_max_14_fsm <= __reduce_max_14_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_24_source_7_source_ram_renable <= 0;
      _stream_conv2d_24_source_7_source_fifo_deq <= 0;
      _stream_conv2d_24_source_7_idle <= 1;
      _stream_conv2d_24_source_9_source_ram_renable <= 0;
      _stream_conv2d_24_source_9_source_fifo_deq <= 0;
      _stream_conv2d_24_source_9_idle <= 1;
      _stream_conv2d_24_source_11_source_ram_renable <= 0;
      _stream_conv2d_24_source_11_source_fifo_deq <= 0;
      _stream_conv2d_24_source_11_idle <= 1;
      _stream_conv2d_24_source_13_source_ram_renable <= 0;
      _stream_conv2d_24_source_13_source_fifo_deq <= 0;
      _stream_conv2d_24_source_13_idle <= 1;
      _stream_conv2d_24_source_15_source_ram_renable <= 0;
      _stream_conv2d_24_source_15_source_fifo_deq <= 0;
      _stream_conv2d_24_source_15_idle <= 1;
      _stream_conv2d_24_source_20_source_ram_renable <= 0;
      _stream_conv2d_24_source_20_source_fifo_deq <= 0;
      _stream_conv2d_24_source_20_idle <= 1;
      _stream_conv2d_24_source_21_source_ram_renable <= 0;
      _stream_conv2d_24_source_21_source_fifo_deq <= 0;
      _stream_conv2d_24_source_21_idle <= 1;
      _stream_conv2d_24_source_22_source_ram_renable <= 0;
      _stream_conv2d_24_source_22_source_fifo_deq <= 0;
      _stream_conv2d_24_source_22_idle <= 1;
      _stream_conv2d_24_source_23_source_ram_renable <= 0;
      _stream_conv2d_24_source_23_source_fifo_deq <= 0;
      _stream_conv2d_24_source_23_idle <= 1;
      _stream_conv2d_24_source_24_source_ram_renable <= 0;
      _stream_conv2d_24_source_24_source_fifo_deq <= 0;
      _stream_conv2d_24_source_24_idle <= 1;
      _stream_conv2d_24_source_25_source_ram_renable <= 0;
      _stream_conv2d_24_source_25_source_fifo_deq <= 0;
      _stream_conv2d_24_source_25_idle <= 1;
      _stream_conv2d_24_source_26_source_ram_renable <= 0;
      _stream_conv2d_24_source_26_source_fifo_deq <= 0;
      _stream_conv2d_24_source_26_idle <= 1;
      _stream_conv2d_24_source_27_source_ram_renable <= 0;
      _stream_conv2d_24_source_27_source_fifo_deq <= 0;
      _stream_conv2d_24_source_27_idle <= 1;
      _stream_conv2d_24_source_28_source_ram_renable <= 0;
      _stream_conv2d_24_source_28_source_fifo_deq <= 0;
      _stream_conv2d_24_source_28_idle <= 1;
      _stream_conv2d_24_source_29_source_ram_renable <= 0;
      _stream_conv2d_24_source_29_source_fifo_deq <= 0;
      _stream_conv2d_24_source_29_idle <= 1;
      _stream_conv2d_24_source_30_source_ram_renable <= 0;
      _stream_conv2d_24_source_30_source_fifo_deq <= 0;
      _stream_conv2d_24_source_30_idle <= 1;
      _stream_conv2d_24_source_31_source_ram_renable <= 0;
      _stream_conv2d_24_source_31_source_fifo_deq <= 0;
      _stream_conv2d_24_source_31_idle <= 1;
      _stream_conv2d_24_source_32_source_ram_renable <= 0;
      _stream_conv2d_24_source_32_source_fifo_deq <= 0;
      _stream_conv2d_24_source_32_idle <= 1;
      _stream_conv2d_24_source_33_source_ram_renable <= 0;
      _stream_conv2d_24_source_33_source_fifo_deq <= 0;
      _stream_conv2d_24_source_33_idle <= 1;
      _stream_conv2d_24_source_34_source_ram_renable <= 0;
      _stream_conv2d_24_source_34_source_fifo_deq <= 0;
      _stream_conv2d_24_source_34_idle <= 1;
      _stream_conv2d_24_source_35_source_ram_renable <= 0;
      _stream_conv2d_24_source_35_source_fifo_deq <= 0;
      _stream_conv2d_24_source_35_idle <= 1;
      _stream_conv2d_24_source_36_source_ram_renable <= 0;
      _stream_conv2d_24_source_36_source_fifo_deq <= 0;
      _stream_conv2d_24_source_36_idle <= 1;
      _stream_conv2d_24_source_37_source_ram_renable <= 0;
      _stream_conv2d_24_source_37_source_fifo_deq <= 0;
      _stream_conv2d_24_source_37_idle <= 1;
      _stream_conv2d_24_sink_50_sink_wenable <= 0;
      _stream_conv2d_24_sink_50_sink_fifo_enq <= 0;
      _stream_conv2d_24_sink_51_sink_wenable <= 0;
      _stream_conv2d_24_sink_51_sink_fifo_enq <= 0;
      __stream_conv2d_24_stream_ivalid_1 <= 0;
      __stream_conv2d_24_stream_ivalid_2 <= 0;
      __stream_conv2d_24_stream_ivalid_3 <= 0;
      __stream_conv2d_24_stream_ivalid_4 <= 0;
      __stream_conv2d_24_stream_ivalid_5 <= 0;
      __stream_conv2d_24_stream_ivalid_6 <= 0;
      __stream_conv2d_24_stream_ivalid_7 <= 0;
      __stream_conv2d_24_stream_ivalid_8 <= 0;
      __stream_conv2d_24_stream_ivalid_9 <= 0;
      __stream_conv2d_24_stream_ivalid_10 <= 0;
      __stream_conv2d_24_stream_ivalid_11 <= 0;
      __stream_conv2d_24_stream_ivalid_12 <= 0;
      __stream_conv2d_24_stream_ivalid_13 <= 0;
      __stream_conv2d_24_stream_ivalid_14 <= 0;
      __stream_conv2d_24_stream_ivalid_15 <= 0;
      __stream_conv2d_24_stream_ivalid_16 <= 0;
      __stream_conv2d_24_stream_ivalid_17 <= 0;
      __stream_conv2d_24_stream_ivalid_18 <= 0;
      __stream_conv2d_24_stream_ivalid_19 <= 0;
      __stream_conv2d_24_stream_ivalid_20 <= 0;
      __stream_conv2d_24_stream_ivalid_21 <= 0;
      __stream_conv2d_24_stream_ivalid_22 <= 0;
      __stream_conv2d_24_stream_ivalid_23 <= 0;
      __stream_conv2d_24_stream_ivalid_24 <= 0;
      __stream_conv2d_24_stream_ivalid_25 <= 0;
      __stream_conv2d_24_stream_ivalid_26 <= 0;
      __stream_conv2d_24_stream_ivalid_27 <= 0;
      __stream_conv2d_24_stream_ivalid_28 <= 0;
      __stream_conv2d_24_stream_ivalid_29 <= 0;
      __stream_conv2d_24_stream_ivalid_30 <= 0;
      __stream_conv2d_24_stream_ivalid_31 <= 0;
      _eq_data_367 <= 0;
      _eq_data_371 <= 0;
      _eq_data_374 <= 0;
      _eq_data_377 <= 0;
      _eq_data_381 <= 0;
      _eq_data_384 <= 0;
      _eq_data_387 <= 0;
      _eq_data_391 <= 0;
      _eq_data_394 <= 0;
      _eq_data_397 <= 0;
      _eq_data_401 <= 0;
      _eq_data_404 <= 0;
      _eq_data_407 <= 0;
      _eq_data_411 <= 0;
      _eq_data_414 <= 0;
      _eq_data_417 <= 0;
      _eq_data_421 <= 0;
      _eq_data_424 <= 0;
      _eq_data_427 <= 0;
      _eq_data_431 <= 0;
      _eq_data_434 <= 0;
      _eq_data_437 <= 0;
      _eq_data_441 <= 0;
      _eq_data_444 <= 0;
      _eq_data_447 <= 0;
      _eq_data_451 <= 0;
      _eq_data_454 <= 0;
      _eq_data_457 <= 0;
      _eq_data_461 <= 0;
      _eq_data_464 <= 0;
      _eq_data_467 <= 0;
      _eq_data_471 <= 0;
      _eq_data_474 <= 0;
      _eq_data_477 <= 0;
      _eq_data_481 <= 0;
      _eq_data_484 <= 0;
      _eq_data_487 <= 0;
      _eq_data_491 <= 0;
      _eq_data_494 <= 0;
      _eq_data_497 <= 0;
      _eq_data_501 <= 0;
      _eq_data_504 <= 0;
      _eq_data_507 <= 0;
      _eq_data_511 <= 0;
      _eq_data_514 <= 0;
      _eq_data_517 <= 0;
      _eq_data_521 <= 0;
      _eq_data_524 <= 0;
      _eq_data_527 <= 0;
      _eq_data_531 <= 0;
      _eq_data_534 <= 0;
      _eq_data_537 <= 0;
      _eq_data_541 <= 0;
      _eq_data_544 <= 0;
      _plus_data_699 <= 0;
      _plus_data_718 <= 0;
      _plus_data_737 <= 0;
      _plus_data_756 <= 0;
      _plus_data_775 <= 0;
      _plus_data_794 <= 0;
      _plus_data_813 <= 0;
      _plus_data_832 <= 0;
      _plus_data_851 <= 0;
      _plus_data_867 <= 0;
      _plus_data_886 <= 0;
      __delay_data_1038__variable_360 <= 0;
      __delay_data_1039__variable_359 <= 0;
      __delay_data_1040__variable_358 <= 0;
      __delay_data_1041__variable_363 <= 0;
      __delay_data_1042__variable_362 <= 0;
      __delay_data_1043__variable_361 <= 0;
      __delay_data_1044__variable_366 <= 0;
      __delay_data_1045__variable_365 <= 0;
      __delay_data_1046__variable_364 <= 0;
      __delay_data_1047_pointer_646 <= 0;
      __delay_data_1048_reinterpretcast_637 <= 0;
      __delay_data_1049_pointer_648 <= 0;
      __delay_data_1050_reinterpretcast_638 <= 0;
      __delay_data_1051_pointer_650 <= 0;
      __delay_data_1052_reinterpretcast_639 <= 0;
      __delay_data_1053_pointer_652 <= 0;
      __delay_data_1054_reinterpretcast_640 <= 0;
      __delay_data_1055_pointer_654 <= 0;
      __delay_data_1056_reinterpretcast_641 <= 0;
      __delay_data_1057_pointer_656 <= 0;
      __delay_data_1058_reinterpretcast_642 <= 0;
      __delay_data_1059_pointer_658 <= 0;
      __delay_data_1060_reinterpretcast_643 <= 0;
      __delay_data_1061_pointer_660 <= 0;
      __delay_data_1062_reinterpretcast_644 <= 0;
      __delay_data_1063_pointer_662 <= 0;
      __delay_data_1064_reinterpretcast_645 <= 0;
      __delay_data_1065__variable_309 <= 0;
      __delay_data_1090__variable_304 <= 0;
      __delay_data_1103_cond_325 <= 0;
      __delay_data_1122_cond_332 <= 0;
      __delay_data_1066__delay_1065__variable_309 <= 0;
      __delay_data_1078_plus_867 <= 0;
      __delay_data_1091__delay_1090__variable_304 <= 0;
      __delay_data_1104__delay_1103_cond_325 <= 0;
      __delay_data_1123__delay_1122_cond_332 <= 0;
      __delay_data_1142_plus_886 <= 0;
      __delay_data_1067__delay_1066__delay_1065__variable_309 <= 0;
      __delay_data_1079__delay_1078_plus_867 <= 0;
      __delay_data_1092__delay_1091__delay_1090__variable_304 <= 0;
      __delay_data_1105__delay_1104__delay_1103_cond_325 <= 0;
      __delay_data_1124__delay_1123__delay_1122_cond_332 <= 0;
      __delay_data_1143__delay_1142_plus_886 <= 0;
      __delay_data_1068__delay_1067__delay_1066____variable_309 <= 0;
      __delay_data_1080__delay_1079__delay_1078_plus_867 <= 0;
      __delay_data_1093__delay_1092__delay_1091____variable_304 <= 0;
      __delay_data_1106__delay_1105__delay_1104__delay_1103_cond_325 <= 0;
      __delay_data_1125__delay_1124__delay_1123__delay_1122_cond_332 <= 0;
      __delay_data_1144__delay_1143__delay_1142_plus_886 <= 0;
      __delay_data_1069__delay_1068__delay_1067____variable_309 <= 0;
      __delay_data_1081__delay_1080__delay_1079__delay_1078_plus_867 <= 0;
      __delay_data_1094__delay_1093__delay_1092____variable_304 <= 0;
      __delay_data_1107__delay_1106__delay_1105__delay_1104___cond_325 <= 0;
      __delay_data_1126__delay_1125__delay_1124__delay_1123___cond_332 <= 0;
      __delay_data_1145__delay_1144__delay_1143__delay_1142_plus_886 <= 0;
      __delay_data_1070__delay_1069__delay_1068____variable_309 <= 0;
      __delay_data_1082__delay_1081__delay_1080__delay_1079___plus_867 <= 0;
      __delay_data_1095__delay_1094__delay_1093____variable_304 <= 0;
      __delay_data_1108__delay_1107__delay_1106__delay_1105___cond_325 <= 0;
      __delay_data_1127__delay_1126__delay_1125__delay_1124___cond_332 <= 0;
      __delay_data_1146__delay_1145__delay_1144__delay_1143___plus_886 <= 0;
      __delay_data_1071__delay_1070__delay_1069____variable_309 <= 0;
      __delay_data_1083__delay_1082__delay_1081__delay_1080___plus_867 <= 0;
      __delay_data_1096__delay_1095__delay_1094____variable_304 <= 0;
      __delay_data_1109__delay_1108__delay_1107__delay_1106___cond_325 <= 0;
      __delay_data_1128__delay_1127__delay_1126__delay_1125___cond_332 <= 0;
      __delay_data_1147__delay_1146__delay_1145__delay_1144___plus_886 <= 0;
      __delay_data_1072__delay_1071__delay_1070____variable_309 <= 0;
      __delay_data_1084__delay_1083__delay_1082__delay_1081___plus_867 <= 0;
      __delay_data_1097__delay_1096__delay_1095____variable_304 <= 0;
      __delay_data_1110__delay_1109__delay_1108__delay_1107___cond_325 <= 0;
      __delay_data_1129__delay_1128__delay_1127__delay_1126___cond_332 <= 0;
      __delay_data_1148__delay_1147__delay_1146__delay_1145___plus_886 <= 0;
      __delay_data_1073__delay_1072__delay_1071____variable_309 <= 0;
      __delay_data_1085__delay_1084__delay_1083__delay_1082___plus_867 <= 0;
      __delay_data_1098__delay_1097__delay_1096____variable_304 <= 0;
      __delay_data_1111__delay_1110__delay_1109__delay_1108___cond_325 <= 0;
      __delay_data_1130__delay_1129__delay_1128__delay_1127___cond_332 <= 0;
      __delay_data_1149__delay_1148__delay_1147__delay_1146___plus_886 <= 0;
      __delay_data_1074__delay_1073__delay_1072____variable_309 <= 0;
      __delay_data_1086__delay_1085__delay_1084__delay_1083___plus_867 <= 0;
      __delay_data_1099__delay_1098__delay_1097____variable_304 <= 0;
      __delay_data_1112__delay_1111__delay_1110__delay_1109___cond_325 <= 0;
      __delay_data_1131__delay_1130__delay_1129__delay_1128___cond_332 <= 0;
      __delay_data_1150__delay_1149__delay_1148__delay_1147___plus_886 <= 0;
      __delay_data_1075__delay_1074__delay_1073____variable_309 <= 0;
      __delay_data_1087__delay_1086__delay_1085__delay_1084___plus_867 <= 0;
      __delay_data_1100__delay_1099__delay_1098____variable_304 <= 0;
      __delay_data_1113__delay_1112__delay_1111__delay_1110___cond_325 <= 0;
      __delay_data_1132__delay_1131__delay_1130__delay_1129___cond_332 <= 0;
      __delay_data_1151__delay_1150__delay_1149__delay_1148___plus_886 <= 0;
      __delay_data_1076__delay_1075__delay_1074____variable_309 <= 0;
      __delay_data_1088__delay_1087__delay_1086__delay_1085___plus_867 <= 0;
      __delay_data_1101__delay_1100__delay_1099____variable_304 <= 0;
      __delay_data_1114__delay_1113__delay_1112__delay_1111___cond_325 <= 0;
      __delay_data_1133__delay_1132__delay_1131__delay_1130___cond_332 <= 0;
      __delay_data_1152__delay_1151__delay_1150__delay_1149___plus_886 <= 0;
      __delay_data_1077__delay_1076__delay_1075____variable_309 <= 0;
      __delay_data_1089__delay_1088__delay_1087__delay_1086___plus_867 <= 0;
      __delay_data_1102__delay_1101__delay_1100____variable_304 <= 0;
      __delay_data_1115__delay_1114__delay_1113__delay_1112___cond_325 <= 0;
      __delay_data_1134__delay_1133__delay_1132__delay_1131___cond_332 <= 0;
      __delay_data_1153__delay_1152__delay_1151__delay_1150___plus_886 <= 0;
      __delay_data_1116__delay_1115__delay_1114__delay_1113___cond_325 <= 0;
      __delay_data_1135__delay_1134__delay_1133__delay_1132___cond_332 <= 0;
      __delay_data_1154__delay_1153__delay_1152__delay_1151___plus_886 <= 0;
      __delay_data_1117__delay_1116__delay_1115__delay_1114___cond_325 <= 0;
      __delay_data_1136__delay_1135__delay_1134__delay_1133___cond_332 <= 0;
      __delay_data_1155__delay_1154__delay_1153__delay_1152___plus_886 <= 0;
      __delay_data_1118__delay_1117__delay_1116__delay_1115___cond_325 <= 0;
      __delay_data_1137__delay_1136__delay_1135__delay_1134___cond_332 <= 0;
      __delay_data_1156__delay_1155__delay_1154__delay_1153___plus_886 <= 0;
      __delay_data_1119__delay_1118__delay_1117__delay_1116___cond_325 <= 0;
      __delay_data_1138__delay_1137__delay_1136__delay_1135___cond_332 <= 0;
      __delay_data_1157__delay_1156__delay_1155__delay_1154___plus_886 <= 0;
      __delay_data_1120__delay_1119__delay_1118__delay_1117___cond_325 <= 0;
      __delay_data_1139__delay_1138__delay_1137__delay_1136___cond_332 <= 0;
      __delay_data_1158__delay_1157__delay_1156__delay_1155___plus_886 <= 0;
      __delay_data_1121__delay_1120__delay_1119__delay_1118___cond_325 <= 0;
      __delay_data_1140__delay_1139__delay_1138__delay_1137___cond_332 <= 0;
      __delay_data_1159__delay_1158__delay_1157__delay_1156___plus_886 <= 0;
      _plus_data_870 <= 0;
      __delay_data_1141__delay_1140__delay_1139__delay_1138___cond_332 <= 0;
      __delay_data_1160__delay_1159__delay_1158__delay_1157___plus_886 <= 0;
      __delay_data_1162__substreamoutput_869 <= 0;
      __delay_data_1163__delay_1162__substreamoutput_869 <= 0;
      __delay_data_1164__delay_1163__delay_1162__substreamoutput_869 <= 0;
      __delay_data_1165__delay_1164__delay_1163____substreamoutput_869 <= 0;
      __delay_data_1166__delay_1165__delay_1164____substreamoutput_869 <= 0;
      __delay_data_1167__delay_1166__delay_1165____substreamoutput_869 <= 0;
      __delay_data_1168__delay_1167__delay_1166____substreamoutput_869 <= 0;
      __delay_data_1169__delay_1168__delay_1167____substreamoutput_869 <= 0;
      __delay_data_1170__delay_1169__delay_1168____substreamoutput_869 <= 0;
      __delay_data_1171__delay_1170__delay_1169____substreamoutput_869 <= 0;
      _greaterthan_data_889 <= 0;
      __delay_data_1161__substreamoutput_887 <= 0;
      __delay_data_1172__delay_1171__delay_1170____substreamoutput_869 <= 0;
      _cond_data_891 <= 0;
      __delay_data_1173__delay_1172__delay_1171____substreamoutput_869 <= 0;
      _stream_conv2d_24_parameter_0_next_parameter_data <= 0;
      __variable_wdata_304 <= 0;
      _stream_conv2d_24_parameter_1_next_parameter_data <= 0;
      __variable_wdata_305 <= 0;
      _stream_conv2d_24_parameter_2_next_parameter_data <= 0;
      __variable_wdata_306 <= 0;
      _stream_conv2d_24_parameter_3_next_parameter_data <= 0;
      __variable_wdata_307 <= 0;
      _stream_conv2d_24_parameter_4_next_parameter_data <= 0;
      __variable_wdata_308 <= 0;
      _stream_conv2d_24_parameter_6_next_parameter_data <= 0;
      __variable_wdata_319 <= 0;
      _stream_conv2d_24_source_7_source_mode <= 5'b0;
      _stream_conv2d_24_source_7_source_offset <= 0;
      _source_stream_conv2d_24_source_7_pat_size_0 <= 0;
      _source_stream_conv2d_24_source_7_pat_stride_0 <= 0;
      _source_stream_conv2d_24_source_7_pat_size_1 <= 0;
      _source_stream_conv2d_24_source_7_pat_stride_1 <= 0;
      _source_stream_conv2d_24_source_7_pat_size_2 <= 0;
      _source_stream_conv2d_24_source_7_pat_stride_2 <= 0;
      _source_stream_conv2d_24_source_7_pat_size_3 <= 0;
      _source_stream_conv2d_24_source_7_pat_stride_3 <= 0;
      _stream_conv2d_24_source_7_source_sel <= 0;
      _stream_conv2d_24_source_7_source_offset_buf <= 0;
      _source_stream_conv2d_24_source_7_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_24_source_7_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_24_source_7_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_24_source_7_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_24_source_7_pat_count_0 <= 0;
      _source_stream_conv2d_24_source_7_pat_count_1 <= 0;
      _source_stream_conv2d_24_source_7_pat_count_2 <= 0;
      _source_stream_conv2d_24_source_7_pat_count_3 <= 0;
      _source_stream_conv2d_24_source_7_pat_size_buf_0 <= 0;
      _source_stream_conv2d_24_source_7_pat_size_buf_1 <= 0;
      _source_stream_conv2d_24_source_7_pat_size_buf_2 <= 0;
      _source_stream_conv2d_24_source_7_pat_size_buf_3 <= 0;
      _source_stream_conv2d_24_source_7_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_24_source_7_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_24_source_7_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_24_source_7_pat_stride_buf_3 <= 0;
      __variable_wdata_320 <= 0;
      _stream_conv2d_24_source_7_source_ram_raddr <= 0;
      _stream_conv2d_24_parameter_8_next_parameter_data <= 0;
      __variable_wdata_326 <= 0;
      _stream_conv2d_24_source_9_source_mode <= 5'b0;
      _stream_conv2d_24_source_9_source_offset <= 0;
      _source_stream_conv2d_24_source_9_pat_size_0 <= 0;
      _source_stream_conv2d_24_source_9_pat_stride_0 <= 0;
      _source_stream_conv2d_24_source_9_pat_size_1 <= 0;
      _source_stream_conv2d_24_source_9_pat_stride_1 <= 0;
      _source_stream_conv2d_24_source_9_pat_size_2 <= 0;
      _source_stream_conv2d_24_source_9_pat_stride_2 <= 0;
      _source_stream_conv2d_24_source_9_pat_size_3 <= 0;
      _source_stream_conv2d_24_source_9_pat_stride_3 <= 0;
      _stream_conv2d_24_source_9_source_sel <= 0;
      _stream_conv2d_24_source_9_source_offset_buf <= 0;
      _source_stream_conv2d_24_source_9_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_24_source_9_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_24_source_9_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_24_source_9_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_24_source_9_pat_count_0 <= 0;
      _source_stream_conv2d_24_source_9_pat_count_1 <= 0;
      _source_stream_conv2d_24_source_9_pat_count_2 <= 0;
      _source_stream_conv2d_24_source_9_pat_count_3 <= 0;
      _source_stream_conv2d_24_source_9_pat_size_buf_0 <= 0;
      _source_stream_conv2d_24_source_9_pat_size_buf_1 <= 0;
      _source_stream_conv2d_24_source_9_pat_size_buf_2 <= 0;
      _source_stream_conv2d_24_source_9_pat_size_buf_3 <= 0;
      _source_stream_conv2d_24_source_9_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_24_source_9_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_24_source_9_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_24_source_9_pat_stride_buf_3 <= 0;
      __variable_wdata_327 <= 0;
      _stream_conv2d_24_source_9_source_ram_raddr <= 0;
      _stream_conv2d_24_parameter_10_next_parameter_data <= 0;
      __variable_wdata_333 <= 0;
      _stream_conv2d_24_source_11_source_mode <= 5'b0;
      _stream_conv2d_24_source_11_source_empty_data <= 0;
      __variable_wdata_334 <= 0;
      _stream_conv2d_24_parameter_12_next_parameter_data <= 0;
      __variable_wdata_340 <= 0;
      _stream_conv2d_24_source_13_source_mode <= 5'b0;
      _stream_conv2d_24_source_13_source_empty_data <= 0;
      __variable_wdata_341 <= 0;
      _stream_conv2d_24_parameter_14_next_parameter_data <= 0;
      __variable_wdata_347 <= 0;
      _stream_conv2d_24_source_15_source_mode <= 5'b0;
      _stream_conv2d_24_source_15_source_empty_data <= 0;
      __variable_wdata_348 <= 0;
      _stream_conv2d_24_parameter_16_next_parameter_data <= 0;
      __variable_wdata_354 <= 0;
      _stream_conv2d_24_parameter_17_next_parameter_data <= 0;
      __variable_wdata_355 <= 0;
      _stream_conv2d_24_parameter_18_next_parameter_data <= 0;
      __variable_wdata_356 <= 0;
      _stream_conv2d_24_parameter_19_next_parameter_data <= 0;
      __variable_wdata_357 <= 0;
      _stream_conv2d_24_source_20_source_mode <= 5'b0;
      _stream_conv2d_24_source_20_source_offset <= 0;
      _source_stream_conv2d_24_source_20_pat_size_0 <= 0;
      _source_stream_conv2d_24_source_20_pat_stride_0 <= 0;
      _source_stream_conv2d_24_source_20_pat_size_1 <= 0;
      _source_stream_conv2d_24_source_20_pat_stride_1 <= 0;
      _source_stream_conv2d_24_source_20_pat_size_2 <= 0;
      _source_stream_conv2d_24_source_20_pat_stride_2 <= 0;
      _source_stream_conv2d_24_source_20_pat_size_3 <= 0;
      _source_stream_conv2d_24_source_20_pat_stride_3 <= 0;
      _stream_conv2d_24_source_20_source_sel <= 0;
      _stream_conv2d_24_source_20_source_offset_buf <= 0;
      _source_stream_conv2d_24_source_20_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_24_source_20_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_24_source_20_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_24_source_20_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_24_source_20_pat_count_0 <= 0;
      _source_stream_conv2d_24_source_20_pat_count_1 <= 0;
      _source_stream_conv2d_24_source_20_pat_count_2 <= 0;
      _source_stream_conv2d_24_source_20_pat_count_3 <= 0;
      _source_stream_conv2d_24_source_20_pat_size_buf_0 <= 0;
      _source_stream_conv2d_24_source_20_pat_size_buf_1 <= 0;
      _source_stream_conv2d_24_source_20_pat_size_buf_2 <= 0;
      _source_stream_conv2d_24_source_20_pat_size_buf_3 <= 0;
      _source_stream_conv2d_24_source_20_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_24_source_20_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_24_source_20_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_24_source_20_pat_stride_buf_3 <= 0;
      __variable_wdata_358 <= 0;
      _stream_conv2d_24_source_20_source_ram_raddr <= 0;
      _stream_conv2d_24_source_21_source_mode <= 5'b0;
      _stream_conv2d_24_source_21_source_offset <= 0;
      _source_stream_conv2d_24_source_21_pat_size_0 <= 0;
      _source_stream_conv2d_24_source_21_pat_stride_0 <= 0;
      _source_stream_conv2d_24_source_21_pat_size_1 <= 0;
      _source_stream_conv2d_24_source_21_pat_stride_1 <= 0;
      _source_stream_conv2d_24_source_21_pat_size_2 <= 0;
      _source_stream_conv2d_24_source_21_pat_stride_2 <= 0;
      _source_stream_conv2d_24_source_21_pat_size_3 <= 0;
      _source_stream_conv2d_24_source_21_pat_stride_3 <= 0;
      _stream_conv2d_24_source_21_source_sel <= 0;
      _stream_conv2d_24_source_21_source_offset_buf <= 0;
      _source_stream_conv2d_24_source_21_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_24_source_21_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_24_source_21_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_24_source_21_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_24_source_21_pat_count_0 <= 0;
      _source_stream_conv2d_24_source_21_pat_count_1 <= 0;
      _source_stream_conv2d_24_source_21_pat_count_2 <= 0;
      _source_stream_conv2d_24_source_21_pat_count_3 <= 0;
      _source_stream_conv2d_24_source_21_pat_size_buf_0 <= 0;
      _source_stream_conv2d_24_source_21_pat_size_buf_1 <= 0;
      _source_stream_conv2d_24_source_21_pat_size_buf_2 <= 0;
      _source_stream_conv2d_24_source_21_pat_size_buf_3 <= 0;
      _source_stream_conv2d_24_source_21_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_24_source_21_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_24_source_21_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_24_source_21_pat_stride_buf_3 <= 0;
      __variable_wdata_359 <= 0;
      _stream_conv2d_24_source_21_source_ram_raddr <= 0;
      _stream_conv2d_24_source_22_source_mode <= 5'b0;
      _stream_conv2d_24_source_22_source_offset <= 0;
      _source_stream_conv2d_24_source_22_pat_size_0 <= 0;
      _source_stream_conv2d_24_source_22_pat_stride_0 <= 0;
      _source_stream_conv2d_24_source_22_pat_size_1 <= 0;
      _source_stream_conv2d_24_source_22_pat_stride_1 <= 0;
      _source_stream_conv2d_24_source_22_pat_size_2 <= 0;
      _source_stream_conv2d_24_source_22_pat_stride_2 <= 0;
      _source_stream_conv2d_24_source_22_pat_size_3 <= 0;
      _source_stream_conv2d_24_source_22_pat_stride_3 <= 0;
      _stream_conv2d_24_source_22_source_sel <= 0;
      _stream_conv2d_24_source_22_source_offset_buf <= 0;
      _source_stream_conv2d_24_source_22_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_24_source_22_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_24_source_22_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_24_source_22_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_24_source_22_pat_count_0 <= 0;
      _source_stream_conv2d_24_source_22_pat_count_1 <= 0;
      _source_stream_conv2d_24_source_22_pat_count_2 <= 0;
      _source_stream_conv2d_24_source_22_pat_count_3 <= 0;
      _source_stream_conv2d_24_source_22_pat_size_buf_0 <= 0;
      _source_stream_conv2d_24_source_22_pat_size_buf_1 <= 0;
      _source_stream_conv2d_24_source_22_pat_size_buf_2 <= 0;
      _source_stream_conv2d_24_source_22_pat_size_buf_3 <= 0;
      _source_stream_conv2d_24_source_22_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_24_source_22_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_24_source_22_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_24_source_22_pat_stride_buf_3 <= 0;
      __variable_wdata_360 <= 0;
      _stream_conv2d_24_source_22_source_ram_raddr <= 0;
      _stream_conv2d_24_source_23_source_mode <= 5'b0;
      _stream_conv2d_24_source_23_source_offset <= 0;
      _source_stream_conv2d_24_source_23_pat_size_0 <= 0;
      _source_stream_conv2d_24_source_23_pat_stride_0 <= 0;
      _source_stream_conv2d_24_source_23_pat_size_1 <= 0;
      _source_stream_conv2d_24_source_23_pat_stride_1 <= 0;
      _source_stream_conv2d_24_source_23_pat_size_2 <= 0;
      _source_stream_conv2d_24_source_23_pat_stride_2 <= 0;
      _source_stream_conv2d_24_source_23_pat_size_3 <= 0;
      _source_stream_conv2d_24_source_23_pat_stride_3 <= 0;
      _stream_conv2d_24_source_23_source_sel <= 0;
      _stream_conv2d_24_source_23_source_offset_buf <= 0;
      _source_stream_conv2d_24_source_23_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_24_source_23_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_24_source_23_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_24_source_23_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_24_source_23_pat_count_0 <= 0;
      _source_stream_conv2d_24_source_23_pat_count_1 <= 0;
      _source_stream_conv2d_24_source_23_pat_count_2 <= 0;
      _source_stream_conv2d_24_source_23_pat_count_3 <= 0;
      _source_stream_conv2d_24_source_23_pat_size_buf_0 <= 0;
      _source_stream_conv2d_24_source_23_pat_size_buf_1 <= 0;
      _source_stream_conv2d_24_source_23_pat_size_buf_2 <= 0;
      _source_stream_conv2d_24_source_23_pat_size_buf_3 <= 0;
      _source_stream_conv2d_24_source_23_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_24_source_23_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_24_source_23_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_24_source_23_pat_stride_buf_3 <= 0;
      __variable_wdata_361 <= 0;
      _stream_conv2d_24_source_23_source_ram_raddr <= 0;
      _stream_conv2d_24_source_24_source_mode <= 5'b0;
      _stream_conv2d_24_source_24_source_offset <= 0;
      _source_stream_conv2d_24_source_24_pat_size_0 <= 0;
      _source_stream_conv2d_24_source_24_pat_stride_0 <= 0;
      _source_stream_conv2d_24_source_24_pat_size_1 <= 0;
      _source_stream_conv2d_24_source_24_pat_stride_1 <= 0;
      _source_stream_conv2d_24_source_24_pat_size_2 <= 0;
      _source_stream_conv2d_24_source_24_pat_stride_2 <= 0;
      _source_stream_conv2d_24_source_24_pat_size_3 <= 0;
      _source_stream_conv2d_24_source_24_pat_stride_3 <= 0;
      _stream_conv2d_24_source_24_source_sel <= 0;
      _stream_conv2d_24_source_24_source_offset_buf <= 0;
      _source_stream_conv2d_24_source_24_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_24_source_24_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_24_source_24_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_24_source_24_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_24_source_24_pat_count_0 <= 0;
      _source_stream_conv2d_24_source_24_pat_count_1 <= 0;
      _source_stream_conv2d_24_source_24_pat_count_2 <= 0;
      _source_stream_conv2d_24_source_24_pat_count_3 <= 0;
      _source_stream_conv2d_24_source_24_pat_size_buf_0 <= 0;
      _source_stream_conv2d_24_source_24_pat_size_buf_1 <= 0;
      _source_stream_conv2d_24_source_24_pat_size_buf_2 <= 0;
      _source_stream_conv2d_24_source_24_pat_size_buf_3 <= 0;
      _source_stream_conv2d_24_source_24_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_24_source_24_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_24_source_24_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_24_source_24_pat_stride_buf_3 <= 0;
      __variable_wdata_362 <= 0;
      _stream_conv2d_24_source_24_source_ram_raddr <= 0;
      _stream_conv2d_24_source_25_source_mode <= 5'b0;
      _stream_conv2d_24_source_25_source_offset <= 0;
      _source_stream_conv2d_24_source_25_pat_size_0 <= 0;
      _source_stream_conv2d_24_source_25_pat_stride_0 <= 0;
      _source_stream_conv2d_24_source_25_pat_size_1 <= 0;
      _source_stream_conv2d_24_source_25_pat_stride_1 <= 0;
      _source_stream_conv2d_24_source_25_pat_size_2 <= 0;
      _source_stream_conv2d_24_source_25_pat_stride_2 <= 0;
      _source_stream_conv2d_24_source_25_pat_size_3 <= 0;
      _source_stream_conv2d_24_source_25_pat_stride_3 <= 0;
      _stream_conv2d_24_source_25_source_sel <= 0;
      _stream_conv2d_24_source_25_source_offset_buf <= 0;
      _source_stream_conv2d_24_source_25_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_24_source_25_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_24_source_25_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_24_source_25_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_24_source_25_pat_count_0 <= 0;
      _source_stream_conv2d_24_source_25_pat_count_1 <= 0;
      _source_stream_conv2d_24_source_25_pat_count_2 <= 0;
      _source_stream_conv2d_24_source_25_pat_count_3 <= 0;
      _source_stream_conv2d_24_source_25_pat_size_buf_0 <= 0;
      _source_stream_conv2d_24_source_25_pat_size_buf_1 <= 0;
      _source_stream_conv2d_24_source_25_pat_size_buf_2 <= 0;
      _source_stream_conv2d_24_source_25_pat_size_buf_3 <= 0;
      _source_stream_conv2d_24_source_25_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_24_source_25_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_24_source_25_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_24_source_25_pat_stride_buf_3 <= 0;
      __variable_wdata_363 <= 0;
      _stream_conv2d_24_source_25_source_ram_raddr <= 0;
      _stream_conv2d_24_source_26_source_mode <= 5'b0;
      _stream_conv2d_24_source_26_source_offset <= 0;
      _source_stream_conv2d_24_source_26_pat_size_0 <= 0;
      _source_stream_conv2d_24_source_26_pat_stride_0 <= 0;
      _source_stream_conv2d_24_source_26_pat_size_1 <= 0;
      _source_stream_conv2d_24_source_26_pat_stride_1 <= 0;
      _source_stream_conv2d_24_source_26_pat_size_2 <= 0;
      _source_stream_conv2d_24_source_26_pat_stride_2 <= 0;
      _source_stream_conv2d_24_source_26_pat_size_3 <= 0;
      _source_stream_conv2d_24_source_26_pat_stride_3 <= 0;
      _stream_conv2d_24_source_26_source_sel <= 0;
      _stream_conv2d_24_source_26_source_offset_buf <= 0;
      _source_stream_conv2d_24_source_26_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_24_source_26_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_24_source_26_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_24_source_26_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_24_source_26_pat_count_0 <= 0;
      _source_stream_conv2d_24_source_26_pat_count_1 <= 0;
      _source_stream_conv2d_24_source_26_pat_count_2 <= 0;
      _source_stream_conv2d_24_source_26_pat_count_3 <= 0;
      _source_stream_conv2d_24_source_26_pat_size_buf_0 <= 0;
      _source_stream_conv2d_24_source_26_pat_size_buf_1 <= 0;
      _source_stream_conv2d_24_source_26_pat_size_buf_2 <= 0;
      _source_stream_conv2d_24_source_26_pat_size_buf_3 <= 0;
      _source_stream_conv2d_24_source_26_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_24_source_26_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_24_source_26_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_24_source_26_pat_stride_buf_3 <= 0;
      __variable_wdata_364 <= 0;
      _stream_conv2d_24_source_26_source_ram_raddr <= 0;
      _stream_conv2d_24_source_27_source_mode <= 5'b0;
      _stream_conv2d_24_source_27_source_offset <= 0;
      _source_stream_conv2d_24_source_27_pat_size_0 <= 0;
      _source_stream_conv2d_24_source_27_pat_stride_0 <= 0;
      _source_stream_conv2d_24_source_27_pat_size_1 <= 0;
      _source_stream_conv2d_24_source_27_pat_stride_1 <= 0;
      _source_stream_conv2d_24_source_27_pat_size_2 <= 0;
      _source_stream_conv2d_24_source_27_pat_stride_2 <= 0;
      _source_stream_conv2d_24_source_27_pat_size_3 <= 0;
      _source_stream_conv2d_24_source_27_pat_stride_3 <= 0;
      _stream_conv2d_24_source_27_source_sel <= 0;
      _stream_conv2d_24_source_27_source_offset_buf <= 0;
      _source_stream_conv2d_24_source_27_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_24_source_27_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_24_source_27_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_24_source_27_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_24_source_27_pat_count_0 <= 0;
      _source_stream_conv2d_24_source_27_pat_count_1 <= 0;
      _source_stream_conv2d_24_source_27_pat_count_2 <= 0;
      _source_stream_conv2d_24_source_27_pat_count_3 <= 0;
      _source_stream_conv2d_24_source_27_pat_size_buf_0 <= 0;
      _source_stream_conv2d_24_source_27_pat_size_buf_1 <= 0;
      _source_stream_conv2d_24_source_27_pat_size_buf_2 <= 0;
      _source_stream_conv2d_24_source_27_pat_size_buf_3 <= 0;
      _source_stream_conv2d_24_source_27_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_24_source_27_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_24_source_27_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_24_source_27_pat_stride_buf_3 <= 0;
      __variable_wdata_365 <= 0;
      _stream_conv2d_24_source_27_source_ram_raddr <= 0;
      _stream_conv2d_24_source_28_source_mode <= 5'b0;
      _stream_conv2d_24_source_28_source_offset <= 0;
      _source_stream_conv2d_24_source_28_pat_size_0 <= 0;
      _source_stream_conv2d_24_source_28_pat_stride_0 <= 0;
      _source_stream_conv2d_24_source_28_pat_size_1 <= 0;
      _source_stream_conv2d_24_source_28_pat_stride_1 <= 0;
      _source_stream_conv2d_24_source_28_pat_size_2 <= 0;
      _source_stream_conv2d_24_source_28_pat_stride_2 <= 0;
      _source_stream_conv2d_24_source_28_pat_size_3 <= 0;
      _source_stream_conv2d_24_source_28_pat_stride_3 <= 0;
      _stream_conv2d_24_source_28_source_sel <= 0;
      _stream_conv2d_24_source_28_source_offset_buf <= 0;
      _source_stream_conv2d_24_source_28_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_24_source_28_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_24_source_28_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_24_source_28_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_24_source_28_pat_count_0 <= 0;
      _source_stream_conv2d_24_source_28_pat_count_1 <= 0;
      _source_stream_conv2d_24_source_28_pat_count_2 <= 0;
      _source_stream_conv2d_24_source_28_pat_count_3 <= 0;
      _source_stream_conv2d_24_source_28_pat_size_buf_0 <= 0;
      _source_stream_conv2d_24_source_28_pat_size_buf_1 <= 0;
      _source_stream_conv2d_24_source_28_pat_size_buf_2 <= 0;
      _source_stream_conv2d_24_source_28_pat_size_buf_3 <= 0;
      _source_stream_conv2d_24_source_28_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_24_source_28_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_24_source_28_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_24_source_28_pat_stride_buf_3 <= 0;
      __variable_wdata_366 <= 0;
      _stream_conv2d_24_source_28_source_ram_raddr <= 0;
      _stream_conv2d_24_source_29_source_mode <= 5'b0;
      _stream_conv2d_24_source_29_source_offset <= 0;
      _source_stream_conv2d_24_source_29_pat_size_0 <= 0;
      _source_stream_conv2d_24_source_29_pat_stride_0 <= 0;
      _source_stream_conv2d_24_source_29_pat_size_1 <= 0;
      _source_stream_conv2d_24_source_29_pat_stride_1 <= 0;
      _source_stream_conv2d_24_source_29_pat_size_2 <= 0;
      _source_stream_conv2d_24_source_29_pat_stride_2 <= 0;
      _source_stream_conv2d_24_source_29_pat_size_3 <= 0;
      _source_stream_conv2d_24_source_29_pat_stride_3 <= 0;
      _stream_conv2d_24_source_29_source_sel <= 0;
      _stream_conv2d_24_source_29_source_offset_buf <= 0;
      _source_stream_conv2d_24_source_29_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_24_source_29_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_24_source_29_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_24_source_29_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_24_source_29_pat_count_0 <= 0;
      _source_stream_conv2d_24_source_29_pat_count_1 <= 0;
      _source_stream_conv2d_24_source_29_pat_count_2 <= 0;
      _source_stream_conv2d_24_source_29_pat_count_3 <= 0;
      _source_stream_conv2d_24_source_29_pat_size_buf_0 <= 0;
      _source_stream_conv2d_24_source_29_pat_size_buf_1 <= 0;
      _source_stream_conv2d_24_source_29_pat_size_buf_2 <= 0;
      _source_stream_conv2d_24_source_29_pat_size_buf_3 <= 0;
      _source_stream_conv2d_24_source_29_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_24_source_29_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_24_source_29_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_24_source_29_pat_stride_buf_3 <= 0;
      __variable_wdata_592 <= 0;
      _stream_conv2d_24_source_29_source_ram_raddr <= 0;
      _stream_conv2d_24_source_30_source_mode <= 5'b0;
      _stream_conv2d_24_source_30_source_offset <= 0;
      _source_stream_conv2d_24_source_30_pat_size_0 <= 0;
      _source_stream_conv2d_24_source_30_pat_stride_0 <= 0;
      _source_stream_conv2d_24_source_30_pat_size_1 <= 0;
      _source_stream_conv2d_24_source_30_pat_stride_1 <= 0;
      _source_stream_conv2d_24_source_30_pat_size_2 <= 0;
      _source_stream_conv2d_24_source_30_pat_stride_2 <= 0;
      _source_stream_conv2d_24_source_30_pat_size_3 <= 0;
      _source_stream_conv2d_24_source_30_pat_stride_3 <= 0;
      _stream_conv2d_24_source_30_source_sel <= 0;
      _stream_conv2d_24_source_30_source_offset_buf <= 0;
      _source_stream_conv2d_24_source_30_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_24_source_30_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_24_source_30_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_24_source_30_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_24_source_30_pat_count_0 <= 0;
      _source_stream_conv2d_24_source_30_pat_count_1 <= 0;
      _source_stream_conv2d_24_source_30_pat_count_2 <= 0;
      _source_stream_conv2d_24_source_30_pat_count_3 <= 0;
      _source_stream_conv2d_24_source_30_pat_size_buf_0 <= 0;
      _source_stream_conv2d_24_source_30_pat_size_buf_1 <= 0;
      _source_stream_conv2d_24_source_30_pat_size_buf_2 <= 0;
      _source_stream_conv2d_24_source_30_pat_size_buf_3 <= 0;
      _source_stream_conv2d_24_source_30_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_24_source_30_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_24_source_30_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_24_source_30_pat_stride_buf_3 <= 0;
      __variable_wdata_593 <= 0;
      _stream_conv2d_24_source_30_source_ram_raddr <= 0;
      _stream_conv2d_24_source_31_source_mode <= 5'b0;
      _stream_conv2d_24_source_31_source_offset <= 0;
      _source_stream_conv2d_24_source_31_pat_size_0 <= 0;
      _source_stream_conv2d_24_source_31_pat_stride_0 <= 0;
      _source_stream_conv2d_24_source_31_pat_size_1 <= 0;
      _source_stream_conv2d_24_source_31_pat_stride_1 <= 0;
      _source_stream_conv2d_24_source_31_pat_size_2 <= 0;
      _source_stream_conv2d_24_source_31_pat_stride_2 <= 0;
      _source_stream_conv2d_24_source_31_pat_size_3 <= 0;
      _source_stream_conv2d_24_source_31_pat_stride_3 <= 0;
      _stream_conv2d_24_source_31_source_sel <= 0;
      _stream_conv2d_24_source_31_source_offset_buf <= 0;
      _source_stream_conv2d_24_source_31_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_24_source_31_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_24_source_31_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_24_source_31_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_24_source_31_pat_count_0 <= 0;
      _source_stream_conv2d_24_source_31_pat_count_1 <= 0;
      _source_stream_conv2d_24_source_31_pat_count_2 <= 0;
      _source_stream_conv2d_24_source_31_pat_count_3 <= 0;
      _source_stream_conv2d_24_source_31_pat_size_buf_0 <= 0;
      _source_stream_conv2d_24_source_31_pat_size_buf_1 <= 0;
      _source_stream_conv2d_24_source_31_pat_size_buf_2 <= 0;
      _source_stream_conv2d_24_source_31_pat_size_buf_3 <= 0;
      _source_stream_conv2d_24_source_31_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_24_source_31_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_24_source_31_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_24_source_31_pat_stride_buf_3 <= 0;
      __variable_wdata_594 <= 0;
      _stream_conv2d_24_source_31_source_ram_raddr <= 0;
      _stream_conv2d_24_source_32_source_mode <= 5'b0;
      _stream_conv2d_24_source_32_source_offset <= 0;
      _source_stream_conv2d_24_source_32_pat_size_0 <= 0;
      _source_stream_conv2d_24_source_32_pat_stride_0 <= 0;
      _source_stream_conv2d_24_source_32_pat_size_1 <= 0;
      _source_stream_conv2d_24_source_32_pat_stride_1 <= 0;
      _source_stream_conv2d_24_source_32_pat_size_2 <= 0;
      _source_stream_conv2d_24_source_32_pat_stride_2 <= 0;
      _source_stream_conv2d_24_source_32_pat_size_3 <= 0;
      _source_stream_conv2d_24_source_32_pat_stride_3 <= 0;
      _stream_conv2d_24_source_32_source_sel <= 0;
      _stream_conv2d_24_source_32_source_offset_buf <= 0;
      _source_stream_conv2d_24_source_32_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_24_source_32_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_24_source_32_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_24_source_32_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_24_source_32_pat_count_0 <= 0;
      _source_stream_conv2d_24_source_32_pat_count_1 <= 0;
      _source_stream_conv2d_24_source_32_pat_count_2 <= 0;
      _source_stream_conv2d_24_source_32_pat_count_3 <= 0;
      _source_stream_conv2d_24_source_32_pat_size_buf_0 <= 0;
      _source_stream_conv2d_24_source_32_pat_size_buf_1 <= 0;
      _source_stream_conv2d_24_source_32_pat_size_buf_2 <= 0;
      _source_stream_conv2d_24_source_32_pat_size_buf_3 <= 0;
      _source_stream_conv2d_24_source_32_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_24_source_32_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_24_source_32_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_24_source_32_pat_stride_buf_3 <= 0;
      __variable_wdata_595 <= 0;
      _stream_conv2d_24_source_32_source_ram_raddr <= 0;
      _stream_conv2d_24_source_33_source_mode <= 5'b0;
      _stream_conv2d_24_source_33_source_offset <= 0;
      _source_stream_conv2d_24_source_33_pat_size_0 <= 0;
      _source_stream_conv2d_24_source_33_pat_stride_0 <= 0;
      _source_stream_conv2d_24_source_33_pat_size_1 <= 0;
      _source_stream_conv2d_24_source_33_pat_stride_1 <= 0;
      _source_stream_conv2d_24_source_33_pat_size_2 <= 0;
      _source_stream_conv2d_24_source_33_pat_stride_2 <= 0;
      _source_stream_conv2d_24_source_33_pat_size_3 <= 0;
      _source_stream_conv2d_24_source_33_pat_stride_3 <= 0;
      _stream_conv2d_24_source_33_source_sel <= 0;
      _stream_conv2d_24_source_33_source_offset_buf <= 0;
      _source_stream_conv2d_24_source_33_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_24_source_33_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_24_source_33_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_24_source_33_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_24_source_33_pat_count_0 <= 0;
      _source_stream_conv2d_24_source_33_pat_count_1 <= 0;
      _source_stream_conv2d_24_source_33_pat_count_2 <= 0;
      _source_stream_conv2d_24_source_33_pat_count_3 <= 0;
      _source_stream_conv2d_24_source_33_pat_size_buf_0 <= 0;
      _source_stream_conv2d_24_source_33_pat_size_buf_1 <= 0;
      _source_stream_conv2d_24_source_33_pat_size_buf_2 <= 0;
      _source_stream_conv2d_24_source_33_pat_size_buf_3 <= 0;
      _source_stream_conv2d_24_source_33_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_24_source_33_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_24_source_33_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_24_source_33_pat_stride_buf_3 <= 0;
      __variable_wdata_596 <= 0;
      _stream_conv2d_24_source_33_source_ram_raddr <= 0;
      _stream_conv2d_24_source_34_source_mode <= 5'b0;
      _stream_conv2d_24_source_34_source_offset <= 0;
      _source_stream_conv2d_24_source_34_pat_size_0 <= 0;
      _source_stream_conv2d_24_source_34_pat_stride_0 <= 0;
      _source_stream_conv2d_24_source_34_pat_size_1 <= 0;
      _source_stream_conv2d_24_source_34_pat_stride_1 <= 0;
      _source_stream_conv2d_24_source_34_pat_size_2 <= 0;
      _source_stream_conv2d_24_source_34_pat_stride_2 <= 0;
      _source_stream_conv2d_24_source_34_pat_size_3 <= 0;
      _source_stream_conv2d_24_source_34_pat_stride_3 <= 0;
      _stream_conv2d_24_source_34_source_sel <= 0;
      _stream_conv2d_24_source_34_source_offset_buf <= 0;
      _source_stream_conv2d_24_source_34_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_24_source_34_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_24_source_34_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_24_source_34_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_24_source_34_pat_count_0 <= 0;
      _source_stream_conv2d_24_source_34_pat_count_1 <= 0;
      _source_stream_conv2d_24_source_34_pat_count_2 <= 0;
      _source_stream_conv2d_24_source_34_pat_count_3 <= 0;
      _source_stream_conv2d_24_source_34_pat_size_buf_0 <= 0;
      _source_stream_conv2d_24_source_34_pat_size_buf_1 <= 0;
      _source_stream_conv2d_24_source_34_pat_size_buf_2 <= 0;
      _source_stream_conv2d_24_source_34_pat_size_buf_3 <= 0;
      _source_stream_conv2d_24_source_34_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_24_source_34_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_24_source_34_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_24_source_34_pat_stride_buf_3 <= 0;
      __variable_wdata_597 <= 0;
      _stream_conv2d_24_source_34_source_ram_raddr <= 0;
      _stream_conv2d_24_source_35_source_mode <= 5'b0;
      _stream_conv2d_24_source_35_source_offset <= 0;
      _source_stream_conv2d_24_source_35_pat_size_0 <= 0;
      _source_stream_conv2d_24_source_35_pat_stride_0 <= 0;
      _source_stream_conv2d_24_source_35_pat_size_1 <= 0;
      _source_stream_conv2d_24_source_35_pat_stride_1 <= 0;
      _source_stream_conv2d_24_source_35_pat_size_2 <= 0;
      _source_stream_conv2d_24_source_35_pat_stride_2 <= 0;
      _source_stream_conv2d_24_source_35_pat_size_3 <= 0;
      _source_stream_conv2d_24_source_35_pat_stride_3 <= 0;
      _stream_conv2d_24_source_35_source_sel <= 0;
      _stream_conv2d_24_source_35_source_offset_buf <= 0;
      _source_stream_conv2d_24_source_35_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_24_source_35_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_24_source_35_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_24_source_35_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_24_source_35_pat_count_0 <= 0;
      _source_stream_conv2d_24_source_35_pat_count_1 <= 0;
      _source_stream_conv2d_24_source_35_pat_count_2 <= 0;
      _source_stream_conv2d_24_source_35_pat_count_3 <= 0;
      _source_stream_conv2d_24_source_35_pat_size_buf_0 <= 0;
      _source_stream_conv2d_24_source_35_pat_size_buf_1 <= 0;
      _source_stream_conv2d_24_source_35_pat_size_buf_2 <= 0;
      _source_stream_conv2d_24_source_35_pat_size_buf_3 <= 0;
      _source_stream_conv2d_24_source_35_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_24_source_35_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_24_source_35_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_24_source_35_pat_stride_buf_3 <= 0;
      __variable_wdata_598 <= 0;
      _stream_conv2d_24_source_35_source_ram_raddr <= 0;
      _stream_conv2d_24_source_36_source_mode <= 5'b0;
      _stream_conv2d_24_source_36_source_offset <= 0;
      _source_stream_conv2d_24_source_36_pat_size_0 <= 0;
      _source_stream_conv2d_24_source_36_pat_stride_0 <= 0;
      _source_stream_conv2d_24_source_36_pat_size_1 <= 0;
      _source_stream_conv2d_24_source_36_pat_stride_1 <= 0;
      _source_stream_conv2d_24_source_36_pat_size_2 <= 0;
      _source_stream_conv2d_24_source_36_pat_stride_2 <= 0;
      _source_stream_conv2d_24_source_36_pat_size_3 <= 0;
      _source_stream_conv2d_24_source_36_pat_stride_3 <= 0;
      _stream_conv2d_24_source_36_source_sel <= 0;
      _stream_conv2d_24_source_36_source_offset_buf <= 0;
      _source_stream_conv2d_24_source_36_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_24_source_36_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_24_source_36_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_24_source_36_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_24_source_36_pat_count_0 <= 0;
      _source_stream_conv2d_24_source_36_pat_count_1 <= 0;
      _source_stream_conv2d_24_source_36_pat_count_2 <= 0;
      _source_stream_conv2d_24_source_36_pat_count_3 <= 0;
      _source_stream_conv2d_24_source_36_pat_size_buf_0 <= 0;
      _source_stream_conv2d_24_source_36_pat_size_buf_1 <= 0;
      _source_stream_conv2d_24_source_36_pat_size_buf_2 <= 0;
      _source_stream_conv2d_24_source_36_pat_size_buf_3 <= 0;
      _source_stream_conv2d_24_source_36_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_24_source_36_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_24_source_36_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_24_source_36_pat_stride_buf_3 <= 0;
      __variable_wdata_599 <= 0;
      _stream_conv2d_24_source_36_source_ram_raddr <= 0;
      _stream_conv2d_24_source_37_source_mode <= 5'b0;
      _stream_conv2d_24_source_37_source_offset <= 0;
      _source_stream_conv2d_24_source_37_pat_size_0 <= 0;
      _source_stream_conv2d_24_source_37_pat_stride_0 <= 0;
      _source_stream_conv2d_24_source_37_pat_size_1 <= 0;
      _source_stream_conv2d_24_source_37_pat_stride_1 <= 0;
      _source_stream_conv2d_24_source_37_pat_size_2 <= 0;
      _source_stream_conv2d_24_source_37_pat_stride_2 <= 0;
      _source_stream_conv2d_24_source_37_pat_size_3 <= 0;
      _source_stream_conv2d_24_source_37_pat_stride_3 <= 0;
      _stream_conv2d_24_source_37_source_sel <= 0;
      _stream_conv2d_24_source_37_source_offset_buf <= 0;
      _source_stream_conv2d_24_source_37_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_24_source_37_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_24_source_37_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_24_source_37_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_24_source_37_pat_count_0 <= 0;
      _source_stream_conv2d_24_source_37_pat_count_1 <= 0;
      _source_stream_conv2d_24_source_37_pat_count_2 <= 0;
      _source_stream_conv2d_24_source_37_pat_count_3 <= 0;
      _source_stream_conv2d_24_source_37_pat_size_buf_0 <= 0;
      _source_stream_conv2d_24_source_37_pat_size_buf_1 <= 0;
      _source_stream_conv2d_24_source_37_pat_size_buf_2 <= 0;
      _source_stream_conv2d_24_source_37_pat_size_buf_3 <= 0;
      _source_stream_conv2d_24_source_37_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_24_source_37_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_24_source_37_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_24_source_37_pat_stride_buf_3 <= 0;
      __variable_wdata_600 <= 0;
      _stream_conv2d_24_source_37_source_ram_raddr <= 0;
      _tmp_665 <= 0;
      _tmp_666 <= 0;
      _tmp_667 <= 0;
      _tmp_668 <= 0;
      _tmp_669 <= 0;
      _tmp_670 <= 0;
      _tmp_671 <= 0;
      _tmp_672 <= 0;
      _tmp_673 <= 0;
      _tmp_674 <= 0;
      _tmp_675 <= 0;
      _tmp_676 <= 0;
      _tmp_677 <= 0;
      _tmp_678 <= 0;
      _tmp_679 <= 0;
      _tmp_680 <= 0;
      _tmp_681 <= 0;
      _tmp_682 <= 0;
      _tmp_683 <= 0;
      _tmp_684 <= 0;
      _tmp_685 <= 0;
      _tmp_686 <= 0;
      _tmp_687 <= 0;
      _tmp_688 <= 0;
      _tmp_689 <= 0;
      _tmp_690 <= 0;
      _tmp_691 <= 0;
      _tmp_692 <= 0;
      _tmp_693 <= 0;
      _tmp_694 <= 0;
      _tmp_695 <= 0;
      _tmp_696 <= 0;
      _tmp_697 <= 0;
      _tmp_700 <= 0;
      _tmp_701 <= 0;
      _tmp_702 <= 0;
      _tmp_703 <= 0;
      _tmp_704 <= 0;
      _tmp_705 <= 0;
      _tmp_706 <= 0;
      _tmp_707 <= 0;
      _tmp_708 <= 0;
      _tmp_709 <= 0;
      _tmp_710 <= 0;
      _tmp_711 <= 0;
      _tmp_712 <= 0;
      _tmp_713 <= 0;
      _tmp_714 <= 0;
      _tmp_715 <= 0;
      _tmp_716 <= 0;
      _tmp_717 <= 0;
      _tmp_718 <= 0;
      _tmp_719 <= 0;
      _tmp_720 <= 0;
      _tmp_721 <= 0;
      _tmp_722 <= 0;
      _tmp_723 <= 0;
      _tmp_724 <= 0;
      _tmp_725 <= 0;
      _tmp_726 <= 0;
      _tmp_727 <= 0;
      _tmp_728 <= 0;
      _tmp_729 <= 0;
      _tmp_730 <= 0;
      _tmp_731 <= 0;
      _tmp_732 <= 0;
      _tmp_733 <= 0;
      _tmp_734 <= 0;
      _tmp_735 <= 0;
      _tmp_736 <= 0;
      _tmp_737 <= 0;
      _tmp_738 <= 0;
      _tmp_739 <= 0;
      _tmp_740 <= 0;
      _tmp_741 <= 0;
      _tmp_742 <= 0;
      _tmp_743 <= 0;
      _tmp_744 <= 0;
      _tmp_745 <= 0;
      _tmp_746 <= 0;
      _tmp_747 <= 0;
      _tmp_748 <= 0;
      _tmp_749 <= 0;
      _tmp_750 <= 0;
      _tmp_751 <= 0;
      _tmp_752 <= 0;
      _tmp_753 <= 0;
      _tmp_754 <= 0;
      _tmp_755 <= 0;
      _tmp_756 <= 0;
      _tmp_757 <= 0;
      _tmp_758 <= 0;
      _tmp_759 <= 0;
      _tmp_760 <= 0;
      _tmp_761 <= 0;
      _tmp_762 <= 0;
      _tmp_763 <= 0;
      _tmp_764 <= 0;
      _tmp_765 <= 0;
      _stream_conv2d_24_sink_50_sink_mode <= 5'b0;
      _stream_conv2d_24_sink_50_sink_offset <= 0;
      _stream_conv2d_24_sink_50_sink_size <= 0;
      _stream_conv2d_24_sink_50_sink_stride <= 0;
      _stream_conv2d_24_sink_50_sink_sel <= 0;
      _stream_conv2d_24_sink_50_sink_offset_buf <= 0;
      _stream_conv2d_24_sink_50_sink_size_buf <= 0;
      _stream_conv2d_24_sink_50_sink_stride_buf <= 0;
      _stream_conv2d_24_sink_50_sink_waddr <= 0;
      _stream_conv2d_24_sink_50_sink_count <= 0;
      _stream_conv2d_24_sink_50_sink_wdata <= 0;
      _tmp_1156 <= 0;
      _tmp_1157 <= 0;
      _tmp_1158 <= 0;
      _tmp_1159 <= 0;
      _tmp_1160 <= 0;
      _tmp_1161 <= 0;
      __variable_wdata_309 <= 0;
      _tmp_1162 <= 0;
      _tmp_1163 <= 0;
      _tmp_1164 <= 0;
      _tmp_1165 <= 0;
      _tmp_1168 <= 0;
      _tmp_1171 <= 0;
      _tmp_1172 <= 0;
      _tmp_1173 <= 0;
      _tmp_1174 <= 0;
      _tmp_1175 <= 0;
      _tmp_1176 <= 0;
      _tmp_1177 <= 0;
      _tmp_1178 <= 0;
      _tmp_1179 <= 0;
      _tmp_1180 <= 0;
      _tmp_1181 <= 0;
      _tmp_1182 <= 0;
      _tmp_1183 <= 0;
      _tmp_1184 <= 0;
      _tmp_1185 <= 0;
      _tmp_1186 <= 0;
      _tmp_1187 <= 0;
      _tmp_1188 <= 0;
      _tmp_1189 <= 0;
      _tmp_1190 <= 0;
      _tmp_1191 <= 0;
      _tmp_1192 <= 0;
      _tmp_1193 <= 0;
      _tmp_1194 <= 0;
      _tmp_1195 <= 0;
      _tmp_1196 <= 0;
      _tmp_1197 <= 0;
      _tmp_1198 <= 0;
      _tmp_1199 <= 0;
      _tmp_1200 <= 0;
      _tmp_1201 <= 0;
      _tmp_1202 <= 0;
      _tmp_1203 <= 0;
      _tmp_1204 <= 0;
      _tmp_1205 <= 0;
      _tmp_1206 <= 0;
      _tmp_1207 <= 0;
      _tmp_1208 <= 0;
      _tmp_1209 <= 0;
      _tmp_1210 <= 0;
      _tmp_1211 <= 0;
      _tmp_1212 <= 0;
      _tmp_1213 <= 0;
      _tmp_1214 <= 0;
      _tmp_1215 <= 0;
      _tmp_1216 <= 0;
      _tmp_1217 <= 0;
      _tmp_1218 <= 0;
      _tmp_1219 <= 0;
      _tmp_1220 <= 0;
      _tmp_1221 <= 0;
      _tmp_1222 <= 0;
      _tmp_1223 <= 0;
      _tmp_1224 <= 0;
      _tmp_1225 <= 0;
      _tmp_1226 <= 0;
      _tmp_1227 <= 0;
      _tmp_1228 <= 0;
      _tmp_1229 <= 0;
      _tmp_1230 <= 0;
      _tmp_1231 <= 0;
      _tmp_1232 <= 0;
      _tmp_1233 <= 0;
      _tmp_1234 <= 0;
      _tmp_1235 <= 0;
      _tmp_1236 <= 0;
      _tmp_1237 <= 0;
      _tmp_1238 <= 0;
      _tmp_1239 <= 0;
      _tmp_1240 <= 0;
      _tmp_1241 <= 0;
      _tmp_1242 <= 0;
      _tmp_1243 <= 0;
      _tmp_1244 <= 0;
      _tmp_1245 <= 0;
      _tmp_1246 <= 0;
      _tmp_1247 <= 0;
      _tmp_1248 <= 0;
      _tmp_1249 <= 0;
      _tmp_1250 <= 0;
      _tmp_1251 <= 0;
      _tmp_1252 <= 0;
      _tmp_1253 <= 0;
      _tmp_1254 <= 0;
      _tmp_1255 <= 0;
      _tmp_1256 <= 0;
      _tmp_1257 <= 0;
      _tmp_1258 <= 0;
      _tmp_1259 <= 0;
      _tmp_1260 <= 0;
      _tmp_1261 <= 0;
      _tmp_1262 <= 0;
      _tmp_1263 <= 0;
      _tmp_1264 <= 0;
      _tmp_1265 <= 0;
      _tmp_1266 <= 0;
      _tmp_1267 <= 0;
      _tmp_1268 <= 0;
      _tmp_1269 <= 0;
      _tmp_1270 <= 0;
      _tmp_1271 <= 0;
      _stream_conv2d_24_busy_reg <= 0;
    end else begin
      if(_stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_7_source_ram_renable <= 0;
        _stream_conv2d_24_source_7_source_fifo_deq <= 0;
      end 
      _stream_conv2d_24_source_7_idle <= _stream_conv2d_24_source_7_idle;
      if(_stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_9_source_ram_renable <= 0;
        _stream_conv2d_24_source_9_source_fifo_deq <= 0;
      end 
      _stream_conv2d_24_source_9_idle <= _stream_conv2d_24_source_9_idle;
      if(_stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_11_source_ram_renable <= 0;
        _stream_conv2d_24_source_11_source_fifo_deq <= 0;
      end 
      _stream_conv2d_24_source_11_idle <= _stream_conv2d_24_source_11_idle;
      if(_stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_13_source_ram_renable <= 0;
        _stream_conv2d_24_source_13_source_fifo_deq <= 0;
      end 
      _stream_conv2d_24_source_13_idle <= _stream_conv2d_24_source_13_idle;
      if(_stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_15_source_ram_renable <= 0;
        _stream_conv2d_24_source_15_source_fifo_deq <= 0;
      end 
      _stream_conv2d_24_source_15_idle <= _stream_conv2d_24_source_15_idle;
      if(_stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_20_source_ram_renable <= 0;
        _stream_conv2d_24_source_20_source_fifo_deq <= 0;
      end 
      _stream_conv2d_24_source_20_idle <= _stream_conv2d_24_source_20_idle;
      if(_stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_21_source_ram_renable <= 0;
        _stream_conv2d_24_source_21_source_fifo_deq <= 0;
      end 
      _stream_conv2d_24_source_21_idle <= _stream_conv2d_24_source_21_idle;
      if(_stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_22_source_ram_renable <= 0;
        _stream_conv2d_24_source_22_source_fifo_deq <= 0;
      end 
      _stream_conv2d_24_source_22_idle <= _stream_conv2d_24_source_22_idle;
      if(_stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_23_source_ram_renable <= 0;
        _stream_conv2d_24_source_23_source_fifo_deq <= 0;
      end 
      _stream_conv2d_24_source_23_idle <= _stream_conv2d_24_source_23_idle;
      if(_stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_24_source_ram_renable <= 0;
        _stream_conv2d_24_source_24_source_fifo_deq <= 0;
      end 
      _stream_conv2d_24_source_24_idle <= _stream_conv2d_24_source_24_idle;
      if(_stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_25_source_ram_renable <= 0;
        _stream_conv2d_24_source_25_source_fifo_deq <= 0;
      end 
      _stream_conv2d_24_source_25_idle <= _stream_conv2d_24_source_25_idle;
      if(_stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_26_source_ram_renable <= 0;
        _stream_conv2d_24_source_26_source_fifo_deq <= 0;
      end 
      _stream_conv2d_24_source_26_idle <= _stream_conv2d_24_source_26_idle;
      if(_stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_27_source_ram_renable <= 0;
        _stream_conv2d_24_source_27_source_fifo_deq <= 0;
      end 
      _stream_conv2d_24_source_27_idle <= _stream_conv2d_24_source_27_idle;
      if(_stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_28_source_ram_renable <= 0;
        _stream_conv2d_24_source_28_source_fifo_deq <= 0;
      end 
      _stream_conv2d_24_source_28_idle <= _stream_conv2d_24_source_28_idle;
      if(_stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_29_source_ram_renable <= 0;
        _stream_conv2d_24_source_29_source_fifo_deq <= 0;
      end 
      _stream_conv2d_24_source_29_idle <= _stream_conv2d_24_source_29_idle;
      if(_stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_30_source_ram_renable <= 0;
        _stream_conv2d_24_source_30_source_fifo_deq <= 0;
      end 
      _stream_conv2d_24_source_30_idle <= _stream_conv2d_24_source_30_idle;
      if(_stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_31_source_ram_renable <= 0;
        _stream_conv2d_24_source_31_source_fifo_deq <= 0;
      end 
      _stream_conv2d_24_source_31_idle <= _stream_conv2d_24_source_31_idle;
      if(_stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_32_source_ram_renable <= 0;
        _stream_conv2d_24_source_32_source_fifo_deq <= 0;
      end 
      _stream_conv2d_24_source_32_idle <= _stream_conv2d_24_source_32_idle;
      if(_stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_33_source_ram_renable <= 0;
        _stream_conv2d_24_source_33_source_fifo_deq <= 0;
      end 
      _stream_conv2d_24_source_33_idle <= _stream_conv2d_24_source_33_idle;
      if(_stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_34_source_ram_renable <= 0;
        _stream_conv2d_24_source_34_source_fifo_deq <= 0;
      end 
      _stream_conv2d_24_source_34_idle <= _stream_conv2d_24_source_34_idle;
      if(_stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_35_source_ram_renable <= 0;
        _stream_conv2d_24_source_35_source_fifo_deq <= 0;
      end 
      _stream_conv2d_24_source_35_idle <= _stream_conv2d_24_source_35_idle;
      if(_stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_36_source_ram_renable <= 0;
        _stream_conv2d_24_source_36_source_fifo_deq <= 0;
      end 
      _stream_conv2d_24_source_36_idle <= _stream_conv2d_24_source_36_idle;
      if(_stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_37_source_ram_renable <= 0;
        _stream_conv2d_24_source_37_source_fifo_deq <= 0;
      end 
      _stream_conv2d_24_source_37_idle <= _stream_conv2d_24_source_37_idle;
      if(_stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_sink_50_sink_wenable <= 0;
        _stream_conv2d_24_sink_50_sink_fifo_enq <= 0;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_sink_51_sink_wenable <= 0;
        _stream_conv2d_24_sink_51_sink_fifo_enq <= 0;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __stream_conv2d_24_stream_ivalid_1 <= _stream_conv2d_24_stream_ivalid;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __stream_conv2d_24_stream_ivalid_2 <= __stream_conv2d_24_stream_ivalid_1;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __stream_conv2d_24_stream_ivalid_3 <= __stream_conv2d_24_stream_ivalid_2;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __stream_conv2d_24_stream_ivalid_4 <= __stream_conv2d_24_stream_ivalid_3;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __stream_conv2d_24_stream_ivalid_5 <= __stream_conv2d_24_stream_ivalid_4;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __stream_conv2d_24_stream_ivalid_6 <= __stream_conv2d_24_stream_ivalid_5;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __stream_conv2d_24_stream_ivalid_7 <= __stream_conv2d_24_stream_ivalid_6;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __stream_conv2d_24_stream_ivalid_8 <= __stream_conv2d_24_stream_ivalid_7;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __stream_conv2d_24_stream_ivalid_9 <= __stream_conv2d_24_stream_ivalid_8;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __stream_conv2d_24_stream_ivalid_10 <= __stream_conv2d_24_stream_ivalid_9;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __stream_conv2d_24_stream_ivalid_11 <= __stream_conv2d_24_stream_ivalid_10;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __stream_conv2d_24_stream_ivalid_12 <= __stream_conv2d_24_stream_ivalid_11;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __stream_conv2d_24_stream_ivalid_13 <= __stream_conv2d_24_stream_ivalid_12;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __stream_conv2d_24_stream_ivalid_14 <= __stream_conv2d_24_stream_ivalid_13;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __stream_conv2d_24_stream_ivalid_15 <= __stream_conv2d_24_stream_ivalid_14;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __stream_conv2d_24_stream_ivalid_16 <= __stream_conv2d_24_stream_ivalid_15;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __stream_conv2d_24_stream_ivalid_17 <= __stream_conv2d_24_stream_ivalid_16;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __stream_conv2d_24_stream_ivalid_18 <= __stream_conv2d_24_stream_ivalid_17;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __stream_conv2d_24_stream_ivalid_19 <= __stream_conv2d_24_stream_ivalid_18;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __stream_conv2d_24_stream_ivalid_20 <= __stream_conv2d_24_stream_ivalid_19;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __stream_conv2d_24_stream_ivalid_21 <= __stream_conv2d_24_stream_ivalid_20;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __stream_conv2d_24_stream_ivalid_22 <= __stream_conv2d_24_stream_ivalid_21;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __stream_conv2d_24_stream_ivalid_23 <= __stream_conv2d_24_stream_ivalid_22;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __stream_conv2d_24_stream_ivalid_24 <= __stream_conv2d_24_stream_ivalid_23;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __stream_conv2d_24_stream_ivalid_25 <= __stream_conv2d_24_stream_ivalid_24;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __stream_conv2d_24_stream_ivalid_26 <= __stream_conv2d_24_stream_ivalid_25;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __stream_conv2d_24_stream_ivalid_27 <= __stream_conv2d_24_stream_ivalid_26;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __stream_conv2d_24_stream_ivalid_28 <= __stream_conv2d_24_stream_ivalid_27;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __stream_conv2d_24_stream_ivalid_29 <= __stream_conv2d_24_stream_ivalid_28;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __stream_conv2d_24_stream_ivalid_30 <= __stream_conv2d_24_stream_ivalid_29;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __stream_conv2d_24_stream_ivalid_31 <= __stream_conv2d_24_stream_ivalid_30;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _eq_data_367 <= stream_conv2d_24_parameter_1_data == 3'sd2;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _eq_data_371 <= stream_conv2d_24_parameter_1_data == 2'sd1;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _eq_data_374 <= stream_conv2d_24_parameter_1_data == 1'sd0;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _eq_data_377 <= stream_conv2d_24_parameter_1_data == 3'sd2;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _eq_data_381 <= stream_conv2d_24_parameter_1_data == 2'sd1;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _eq_data_384 <= stream_conv2d_24_parameter_1_data == 1'sd0;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _eq_data_387 <= stream_conv2d_24_parameter_1_data == 3'sd2;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _eq_data_391 <= stream_conv2d_24_parameter_1_data == 2'sd1;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _eq_data_394 <= stream_conv2d_24_parameter_1_data == 1'sd0;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _eq_data_397 <= stream_conv2d_24_parameter_1_data == 3'sd2;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _eq_data_401 <= stream_conv2d_24_parameter_1_data == 2'sd1;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _eq_data_404 <= stream_conv2d_24_parameter_1_data == 1'sd0;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _eq_data_407 <= stream_conv2d_24_parameter_1_data == 3'sd2;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _eq_data_411 <= stream_conv2d_24_parameter_1_data == 2'sd1;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _eq_data_414 <= stream_conv2d_24_parameter_1_data == 1'sd0;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _eq_data_417 <= stream_conv2d_24_parameter_1_data == 3'sd2;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _eq_data_421 <= stream_conv2d_24_parameter_1_data == 2'sd1;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _eq_data_424 <= stream_conv2d_24_parameter_1_data == 1'sd0;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _eq_data_427 <= stream_conv2d_24_parameter_1_data == 3'sd2;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _eq_data_431 <= stream_conv2d_24_parameter_1_data == 2'sd1;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _eq_data_434 <= stream_conv2d_24_parameter_1_data == 1'sd0;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _eq_data_437 <= stream_conv2d_24_parameter_1_data == 3'sd2;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _eq_data_441 <= stream_conv2d_24_parameter_1_data == 2'sd1;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _eq_data_444 <= stream_conv2d_24_parameter_1_data == 1'sd0;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _eq_data_447 <= stream_conv2d_24_parameter_1_data == 3'sd2;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _eq_data_451 <= stream_conv2d_24_parameter_1_data == 2'sd1;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _eq_data_454 <= stream_conv2d_24_parameter_1_data == 1'sd0;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _eq_data_457 <= stream_conv2d_24_parameter_2_data == 3'sd2;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _eq_data_461 <= stream_conv2d_24_parameter_2_data == 2'sd1;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _eq_data_464 <= stream_conv2d_24_parameter_2_data == 1'sd0;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _eq_data_467 <= stream_conv2d_24_parameter_2_data == 3'sd2;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _eq_data_471 <= stream_conv2d_24_parameter_2_data == 2'sd1;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _eq_data_474 <= stream_conv2d_24_parameter_2_data == 1'sd0;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _eq_data_477 <= stream_conv2d_24_parameter_2_data == 3'sd2;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _eq_data_481 <= stream_conv2d_24_parameter_2_data == 2'sd1;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _eq_data_484 <= stream_conv2d_24_parameter_2_data == 1'sd0;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _eq_data_487 <= stream_conv2d_24_parameter_2_data == 3'sd2;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _eq_data_491 <= stream_conv2d_24_parameter_2_data == 2'sd1;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _eq_data_494 <= stream_conv2d_24_parameter_2_data == 1'sd0;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _eq_data_497 <= stream_conv2d_24_parameter_2_data == 3'sd2;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _eq_data_501 <= stream_conv2d_24_parameter_2_data == 2'sd1;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _eq_data_504 <= stream_conv2d_24_parameter_2_data == 1'sd0;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _eq_data_507 <= stream_conv2d_24_parameter_2_data == 3'sd2;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _eq_data_511 <= stream_conv2d_24_parameter_2_data == 2'sd1;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _eq_data_514 <= stream_conv2d_24_parameter_2_data == 1'sd0;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _eq_data_517 <= stream_conv2d_24_parameter_2_data == 3'sd2;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _eq_data_521 <= stream_conv2d_24_parameter_2_data == 2'sd1;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _eq_data_524 <= stream_conv2d_24_parameter_2_data == 1'sd0;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _eq_data_527 <= stream_conv2d_24_parameter_2_data == 3'sd2;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _eq_data_531 <= stream_conv2d_24_parameter_2_data == 2'sd1;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _eq_data_534 <= stream_conv2d_24_parameter_2_data == 1'sd0;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _eq_data_537 <= stream_conv2d_24_parameter_2_data == 3'sd2;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _eq_data_541 <= stream_conv2d_24_parameter_2_data == 2'sd1;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _eq_data_544 <= stream_conv2d_24_parameter_2_data == 1'sd0;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _plus_data_699 <= _cond_data_339 + stream_conv2d_24_parameter_16_data;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _plus_data_718 <= _cond_data_339 + stream_conv2d_24_parameter_16_data;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _plus_data_737 <= _cond_data_339 + stream_conv2d_24_parameter_16_data;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _plus_data_756 <= _cond_data_339 + stream_conv2d_24_parameter_16_data;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _plus_data_775 <= _cond_data_339 + stream_conv2d_24_parameter_16_data;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _plus_data_794 <= _cond_data_339 + stream_conv2d_24_parameter_16_data;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _plus_data_813 <= _cond_data_339 + stream_conv2d_24_parameter_16_data;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _plus_data_832 <= _cond_data_339 + stream_conv2d_24_parameter_16_data;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _plus_data_851 <= _cond_data_339 + stream_conv2d_24_parameter_16_data;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _plus_data_867 <= _cond_data_346 + stream_conv2d_24_parameter_17_data;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _plus_data_886 <= _cond_data_353 + stream_conv2d_24_parameter_18_data;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1038__variable_360 <= stream_conv2d_24_source_22_data;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1039__variable_359 <= stream_conv2d_24_source_21_data;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1040__variable_358 <= stream_conv2d_24_source_20_data;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1041__variable_363 <= stream_conv2d_24_source_25_data;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1042__variable_362 <= stream_conv2d_24_source_24_data;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1043__variable_361 <= stream_conv2d_24_source_23_data;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1044__variable_366 <= stream_conv2d_24_source_28_data;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1045__variable_365 <= stream_conv2d_24_source_27_data;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1046__variable_364 <= stream_conv2d_24_source_26_data;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1047_pointer_646 <= _pointer_data_646;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1048_reinterpretcast_637 <= _reinterpretcast_data_637;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1049_pointer_648 <= _pointer_data_648;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1050_reinterpretcast_638 <= _reinterpretcast_data_638;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1051_pointer_650 <= _pointer_data_650;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1052_reinterpretcast_639 <= _reinterpretcast_data_639;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1053_pointer_652 <= _pointer_data_652;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1054_reinterpretcast_640 <= _reinterpretcast_data_640;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1055_pointer_654 <= _pointer_data_654;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1056_reinterpretcast_641 <= _reinterpretcast_data_641;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1057_pointer_656 <= _pointer_data_656;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1058_reinterpretcast_642 <= _reinterpretcast_data_642;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1059_pointer_658 <= _pointer_data_658;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1060_reinterpretcast_643 <= _reinterpretcast_data_643;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1061_pointer_660 <= _pointer_data_660;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1062_reinterpretcast_644 <= _reinterpretcast_data_644;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1063_pointer_662 <= _pointer_data_662;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1064_reinterpretcast_645 <= _reinterpretcast_data_645;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1065__variable_309 <= stream_conv2d_24__reduce_reset_data;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1090__variable_304 <= stream_conv2d_24_parameter_0_data;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1103_cond_325 <= _cond_data_325;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1122_cond_332 <= _cond_data_332;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1066__delay_1065__variable_309 <= __delay_data_1065__variable_309;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1078_plus_867 <= _plus_data_867;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1091__delay_1090__variable_304 <= __delay_data_1090__variable_304;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1104__delay_1103_cond_325 <= __delay_data_1103_cond_325;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1123__delay_1122_cond_332 <= __delay_data_1122_cond_332;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1142_plus_886 <= _plus_data_886;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1067__delay_1066__delay_1065__variable_309 <= __delay_data_1066__delay_1065__variable_309;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1079__delay_1078_plus_867 <= __delay_data_1078_plus_867;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1092__delay_1091__delay_1090__variable_304 <= __delay_data_1091__delay_1090__variable_304;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1105__delay_1104__delay_1103_cond_325 <= __delay_data_1104__delay_1103_cond_325;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1124__delay_1123__delay_1122_cond_332 <= __delay_data_1123__delay_1122_cond_332;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1143__delay_1142_plus_886 <= __delay_data_1142_plus_886;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1068__delay_1067__delay_1066____variable_309 <= __delay_data_1067__delay_1066__delay_1065__variable_309;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1080__delay_1079__delay_1078_plus_867 <= __delay_data_1079__delay_1078_plus_867;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1093__delay_1092__delay_1091____variable_304 <= __delay_data_1092__delay_1091__delay_1090__variable_304;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1106__delay_1105__delay_1104__delay_1103_cond_325 <= __delay_data_1105__delay_1104__delay_1103_cond_325;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1125__delay_1124__delay_1123__delay_1122_cond_332 <= __delay_data_1124__delay_1123__delay_1122_cond_332;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1144__delay_1143__delay_1142_plus_886 <= __delay_data_1143__delay_1142_plus_886;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1069__delay_1068__delay_1067____variable_309 <= __delay_data_1068__delay_1067__delay_1066____variable_309;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1081__delay_1080__delay_1079__delay_1078_plus_867 <= __delay_data_1080__delay_1079__delay_1078_plus_867;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1094__delay_1093__delay_1092____variable_304 <= __delay_data_1093__delay_1092__delay_1091____variable_304;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1107__delay_1106__delay_1105__delay_1104___cond_325 <= __delay_data_1106__delay_1105__delay_1104__delay_1103_cond_325;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1126__delay_1125__delay_1124__delay_1123___cond_332 <= __delay_data_1125__delay_1124__delay_1123__delay_1122_cond_332;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1145__delay_1144__delay_1143__delay_1142_plus_886 <= __delay_data_1144__delay_1143__delay_1142_plus_886;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1070__delay_1069__delay_1068____variable_309 <= __delay_data_1069__delay_1068__delay_1067____variable_309;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1082__delay_1081__delay_1080__delay_1079___plus_867 <= __delay_data_1081__delay_1080__delay_1079__delay_1078_plus_867;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1095__delay_1094__delay_1093____variable_304 <= __delay_data_1094__delay_1093__delay_1092____variable_304;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1108__delay_1107__delay_1106__delay_1105___cond_325 <= __delay_data_1107__delay_1106__delay_1105__delay_1104___cond_325;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1127__delay_1126__delay_1125__delay_1124___cond_332 <= __delay_data_1126__delay_1125__delay_1124__delay_1123___cond_332;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1146__delay_1145__delay_1144__delay_1143___plus_886 <= __delay_data_1145__delay_1144__delay_1143__delay_1142_plus_886;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1071__delay_1070__delay_1069____variable_309 <= __delay_data_1070__delay_1069__delay_1068____variable_309;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1083__delay_1082__delay_1081__delay_1080___plus_867 <= __delay_data_1082__delay_1081__delay_1080__delay_1079___plus_867;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1096__delay_1095__delay_1094____variable_304 <= __delay_data_1095__delay_1094__delay_1093____variable_304;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1109__delay_1108__delay_1107__delay_1106___cond_325 <= __delay_data_1108__delay_1107__delay_1106__delay_1105___cond_325;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1128__delay_1127__delay_1126__delay_1125___cond_332 <= __delay_data_1127__delay_1126__delay_1125__delay_1124___cond_332;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1147__delay_1146__delay_1145__delay_1144___plus_886 <= __delay_data_1146__delay_1145__delay_1144__delay_1143___plus_886;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1072__delay_1071__delay_1070____variable_309 <= __delay_data_1071__delay_1070__delay_1069____variable_309;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1084__delay_1083__delay_1082__delay_1081___plus_867 <= __delay_data_1083__delay_1082__delay_1081__delay_1080___plus_867;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1097__delay_1096__delay_1095____variable_304 <= __delay_data_1096__delay_1095__delay_1094____variable_304;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1110__delay_1109__delay_1108__delay_1107___cond_325 <= __delay_data_1109__delay_1108__delay_1107__delay_1106___cond_325;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1129__delay_1128__delay_1127__delay_1126___cond_332 <= __delay_data_1128__delay_1127__delay_1126__delay_1125___cond_332;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1148__delay_1147__delay_1146__delay_1145___plus_886 <= __delay_data_1147__delay_1146__delay_1145__delay_1144___plus_886;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1073__delay_1072__delay_1071____variable_309 <= __delay_data_1072__delay_1071__delay_1070____variable_309;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1085__delay_1084__delay_1083__delay_1082___plus_867 <= __delay_data_1084__delay_1083__delay_1082__delay_1081___plus_867;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1098__delay_1097__delay_1096____variable_304 <= __delay_data_1097__delay_1096__delay_1095____variable_304;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1111__delay_1110__delay_1109__delay_1108___cond_325 <= __delay_data_1110__delay_1109__delay_1108__delay_1107___cond_325;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1130__delay_1129__delay_1128__delay_1127___cond_332 <= __delay_data_1129__delay_1128__delay_1127__delay_1126___cond_332;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1149__delay_1148__delay_1147__delay_1146___plus_886 <= __delay_data_1148__delay_1147__delay_1146__delay_1145___plus_886;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1074__delay_1073__delay_1072____variable_309 <= __delay_data_1073__delay_1072__delay_1071____variable_309;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1086__delay_1085__delay_1084__delay_1083___plus_867 <= __delay_data_1085__delay_1084__delay_1083__delay_1082___plus_867;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1099__delay_1098__delay_1097____variable_304 <= __delay_data_1098__delay_1097__delay_1096____variable_304;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1112__delay_1111__delay_1110__delay_1109___cond_325 <= __delay_data_1111__delay_1110__delay_1109__delay_1108___cond_325;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1131__delay_1130__delay_1129__delay_1128___cond_332 <= __delay_data_1130__delay_1129__delay_1128__delay_1127___cond_332;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1150__delay_1149__delay_1148__delay_1147___plus_886 <= __delay_data_1149__delay_1148__delay_1147__delay_1146___plus_886;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1075__delay_1074__delay_1073____variable_309 <= __delay_data_1074__delay_1073__delay_1072____variable_309;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1087__delay_1086__delay_1085__delay_1084___plus_867 <= __delay_data_1086__delay_1085__delay_1084__delay_1083___plus_867;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1100__delay_1099__delay_1098____variable_304 <= __delay_data_1099__delay_1098__delay_1097____variable_304;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1113__delay_1112__delay_1111__delay_1110___cond_325 <= __delay_data_1112__delay_1111__delay_1110__delay_1109___cond_325;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1132__delay_1131__delay_1130__delay_1129___cond_332 <= __delay_data_1131__delay_1130__delay_1129__delay_1128___cond_332;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1151__delay_1150__delay_1149__delay_1148___plus_886 <= __delay_data_1150__delay_1149__delay_1148__delay_1147___plus_886;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1076__delay_1075__delay_1074____variable_309 <= __delay_data_1075__delay_1074__delay_1073____variable_309;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1088__delay_1087__delay_1086__delay_1085___plus_867 <= __delay_data_1087__delay_1086__delay_1085__delay_1084___plus_867;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1101__delay_1100__delay_1099____variable_304 <= __delay_data_1100__delay_1099__delay_1098____variable_304;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1114__delay_1113__delay_1112__delay_1111___cond_325 <= __delay_data_1113__delay_1112__delay_1111__delay_1110___cond_325;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1133__delay_1132__delay_1131__delay_1130___cond_332 <= __delay_data_1132__delay_1131__delay_1130__delay_1129___cond_332;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1152__delay_1151__delay_1150__delay_1149___plus_886 <= __delay_data_1151__delay_1150__delay_1149__delay_1148___plus_886;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1077__delay_1076__delay_1075____variable_309 <= __delay_data_1076__delay_1075__delay_1074____variable_309;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1089__delay_1088__delay_1087__delay_1086___plus_867 <= __delay_data_1088__delay_1087__delay_1086__delay_1085___plus_867;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1102__delay_1101__delay_1100____variable_304 <= __delay_data_1101__delay_1100__delay_1099____variable_304;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1115__delay_1114__delay_1113__delay_1112___cond_325 <= __delay_data_1114__delay_1113__delay_1112__delay_1111___cond_325;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1134__delay_1133__delay_1132__delay_1131___cond_332 <= __delay_data_1133__delay_1132__delay_1131__delay_1130___cond_332;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1153__delay_1152__delay_1151__delay_1150___plus_886 <= __delay_data_1152__delay_1151__delay_1150__delay_1149___plus_886;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1116__delay_1115__delay_1114__delay_1113___cond_325 <= __delay_data_1115__delay_1114__delay_1113__delay_1112___cond_325;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1135__delay_1134__delay_1133__delay_1132___cond_332 <= __delay_data_1134__delay_1133__delay_1132__delay_1131___cond_332;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1154__delay_1153__delay_1152__delay_1151___plus_886 <= __delay_data_1153__delay_1152__delay_1151__delay_1150___plus_886;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1117__delay_1116__delay_1115__delay_1114___cond_325 <= __delay_data_1116__delay_1115__delay_1114__delay_1113___cond_325;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1136__delay_1135__delay_1134__delay_1133___cond_332 <= __delay_data_1135__delay_1134__delay_1133__delay_1132___cond_332;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1155__delay_1154__delay_1153__delay_1152___plus_886 <= __delay_data_1154__delay_1153__delay_1152__delay_1151___plus_886;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1118__delay_1117__delay_1116__delay_1115___cond_325 <= __delay_data_1117__delay_1116__delay_1115__delay_1114___cond_325;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1137__delay_1136__delay_1135__delay_1134___cond_332 <= __delay_data_1136__delay_1135__delay_1134__delay_1133___cond_332;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1156__delay_1155__delay_1154__delay_1153___plus_886 <= __delay_data_1155__delay_1154__delay_1153__delay_1152___plus_886;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1119__delay_1118__delay_1117__delay_1116___cond_325 <= __delay_data_1118__delay_1117__delay_1116__delay_1115___cond_325;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1138__delay_1137__delay_1136__delay_1135___cond_332 <= __delay_data_1137__delay_1136__delay_1135__delay_1134___cond_332;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1157__delay_1156__delay_1155__delay_1154___plus_886 <= __delay_data_1156__delay_1155__delay_1154__delay_1153___plus_886;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1120__delay_1119__delay_1118__delay_1117___cond_325 <= __delay_data_1119__delay_1118__delay_1117__delay_1116___cond_325;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1139__delay_1138__delay_1137__delay_1136___cond_332 <= __delay_data_1138__delay_1137__delay_1136__delay_1135___cond_332;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1158__delay_1157__delay_1156__delay_1155___plus_886 <= __delay_data_1157__delay_1156__delay_1155__delay_1154___plus_886;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1121__delay_1120__delay_1119__delay_1118___cond_325 <= __delay_data_1120__delay_1119__delay_1118__delay_1117___cond_325;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1140__delay_1139__delay_1138__delay_1137___cond_332 <= __delay_data_1139__delay_1138__delay_1137__delay_1136___cond_332;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1159__delay_1158__delay_1157__delay_1156___plus_886 <= __delay_data_1158__delay_1157__delay_1156__delay_1155___plus_886;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _plus_data_870 <= __substreamoutput_data_868 + __delay_data_1121__delay_1120__delay_1119__delay_1118___cond_325;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1141__delay_1140__delay_1139__delay_1138___cond_332 <= __delay_data_1140__delay_1139__delay_1138__delay_1137___cond_332;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1160__delay_1159__delay_1158__delay_1157___plus_886 <= __delay_data_1159__delay_1158__delay_1157__delay_1156___plus_886;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1162__substreamoutput_869 <= __substreamoutput_data_869;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1163__delay_1162__substreamoutput_869 <= __delay_data_1162__substreamoutput_869;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1164__delay_1163__delay_1162__substreamoutput_869 <= __delay_data_1163__delay_1162__substreamoutput_869;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1165__delay_1164__delay_1163____substreamoutput_869 <= __delay_data_1164__delay_1163__delay_1162__substreamoutput_869;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1166__delay_1165__delay_1164____substreamoutput_869 <= __delay_data_1165__delay_1164__delay_1163____substreamoutput_869;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1167__delay_1166__delay_1165____substreamoutput_869 <= __delay_data_1166__delay_1165__delay_1164____substreamoutput_869;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1168__delay_1167__delay_1166____substreamoutput_869 <= __delay_data_1167__delay_1166__delay_1165____substreamoutput_869;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1169__delay_1168__delay_1167____substreamoutput_869 <= __delay_data_1168__delay_1167__delay_1166____substreamoutput_869;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1170__delay_1169__delay_1168____substreamoutput_869 <= __delay_data_1169__delay_1168__delay_1167____substreamoutput_869;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1171__delay_1170__delay_1169____substreamoutput_869 <= __delay_data_1170__delay_1169__delay_1168____substreamoutput_869;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _greaterthan_data_889 <= __substreamoutput_data_887 > 1'sd0;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1161__substreamoutput_887 <= __substreamoutput_data_887;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1172__delay_1171__delay_1170____substreamoutput_869 <= __delay_data_1171__delay_1170__delay_1169____substreamoutput_869;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _cond_data_891 <= (_greaterthan_data_889)? __delay_data_1161__substreamoutput_887 : 1'sd0;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        __delay_data_1173__delay_1172__delay_1171____substreamoutput_869 <= __delay_data_1172__delay_1171__delay_1170____substreamoutput_869;
      end 
      if(_set_flag_397) begin
        _stream_conv2d_24_parameter_0_next_parameter_data <= cparam_conv2d_24_stream_reduce_size;
      end 
      if(_stream_conv2d_24_source_start) begin
        __variable_wdata_304 <= _stream_conv2d_24_parameter_0_next_parameter_data;
      end 
      if(_set_flag_398) begin
        _stream_conv2d_24_parameter_1_next_parameter_data <= conv2d_24_col_select;
      end 
      if(_stream_conv2d_24_source_start) begin
        __variable_wdata_305 <= _stream_conv2d_24_parameter_1_next_parameter_data;
      end 
      if(_set_flag_399) begin
        _stream_conv2d_24_parameter_2_next_parameter_data <= conv2d_24_row_select_buf;
      end 
      if(_stream_conv2d_24_source_start) begin
        __variable_wdata_306 <= _stream_conv2d_24_parameter_2_next_parameter_data;
      end 
      if(_set_flag_400) begin
        _stream_conv2d_24_parameter_3_next_parameter_data <= conv2d_24_stream_pad_masks;
      end 
      if(_stream_conv2d_24_source_start) begin
        __variable_wdata_307 <= _stream_conv2d_24_parameter_3_next_parameter_data;
      end 
      if(_set_flag_401) begin
        _stream_conv2d_24_parameter_4_next_parameter_data <= cparam_conv2d_24_stream_omit_mask;
      end 
      if(_stream_conv2d_24_source_start) begin
        __variable_wdata_308 <= _stream_conv2d_24_parameter_4_next_parameter_data;
      end 
      if(_set_flag_402) begin
        _stream_conv2d_24_parameter_6_next_parameter_data <= cparam_conv2d_24_bias_scala;
      end 
      if(_stream_conv2d_24_source_start) begin
        __variable_wdata_319 <= _stream_conv2d_24_parameter_6_next_parameter_data;
      end 
      if(_set_flag_403) begin
        _stream_conv2d_24_source_7_source_mode <= 5'b10;
        _stream_conv2d_24_source_7_source_offset <= (cparam_conv2d_24_bias_num == 1)? 0 : conv2d_24_och_count_buf;
      end 
      if(_set_flag_403) begin
        _source_stream_conv2d_24_source_7_pat_size_0 <= cparam_conv2d_24_stream_reduce_size;
        _source_stream_conv2d_24_source_7_pat_stride_0 <= 0;
      end 
      if(_set_flag_403) begin
        _source_stream_conv2d_24_source_7_pat_size_1 <= conv2d_24_next_stream_num_ops;
        _source_stream_conv2d_24_source_7_pat_stride_1 <= (cparam_conv2d_24_bias_num == 1)? 0 : 1;
      end 
      if(_set_flag_403) begin
        _source_stream_conv2d_24_source_7_pat_size_2 <= 1;
        _source_stream_conv2d_24_source_7_pat_stride_2 <= 0;
      end 
      if(_set_flag_403) begin
        _source_stream_conv2d_24_source_7_pat_size_3 <= 1;
        _source_stream_conv2d_24_source_7_pat_stride_3 <= 0;
      end 
      if(_set_flag_403) begin
        _stream_conv2d_24_source_7_source_sel <= 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_7_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_7_source_offset_buf <= _stream_conv2d_24_source_7_source_offset;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_7_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_7_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_7_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_7_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_7_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_7_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_7_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_7_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_7_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_7_pat_count_0 <= _source_stream_conv2d_24_source_7_pat_size_0 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_7_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_7_pat_count_1 <= _source_stream_conv2d_24_source_7_pat_size_1 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_7_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_7_pat_count_2 <= _source_stream_conv2d_24_source_7_pat_size_2 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_7_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_7_pat_count_3 <= _source_stream_conv2d_24_source_7_pat_size_3 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_7_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_7_pat_size_buf_0 <= _source_stream_conv2d_24_source_7_pat_size_0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_7_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_7_pat_size_buf_1 <= _source_stream_conv2d_24_source_7_pat_size_1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_7_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_7_pat_size_buf_2 <= _source_stream_conv2d_24_source_7_pat_size_2;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_7_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_7_pat_size_buf_3 <= _source_stream_conv2d_24_source_7_pat_size_3;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_7_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_7_pat_stride_buf_0 <= _source_stream_conv2d_24_source_7_pat_stride_0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_7_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_7_pat_stride_buf_1 <= _source_stream_conv2d_24_source_7_pat_stride_1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_7_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_7_pat_stride_buf_2 <= _source_stream_conv2d_24_source_7_pat_stride_2;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_7_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_7_pat_stride_buf_3 <= _source_stream_conv2d_24_source_7_pat_stride_3;
      end 
      if(_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_busy && _stream_conv2d_24_is_root) begin
        __variable_wdata_320 <= _stream_conv2d_24_source_7_source_ram_rdata;
      end 
      if((_stream_conv2d_24_source_7_source_pat_fsm_0 == 1) && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_7_idle <= 0;
        _stream_conv2d_24_source_7_source_ram_raddr <= _stream_conv2d_24_source_7_source_pat_all_offset;
        _stream_conv2d_24_source_7_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_24_source_7_source_pat_fsm_0 == 1) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_7_pat_cur_offset_0 <= _source_stream_conv2d_24_source_7_pat_cur_offset_0 + _source_stream_conv2d_24_source_7_pat_stride_buf_0;
        _source_stream_conv2d_24_source_7_pat_count_0 <= _source_stream_conv2d_24_source_7_pat_count_0 - 1;
      end 
      if((_stream_conv2d_24_source_7_source_pat_fsm_0 == 1) && (_source_stream_conv2d_24_source_7_pat_count_0 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_7_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_24_source_7_pat_count_0 <= _source_stream_conv2d_24_source_7_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_24_source_7_source_pat_fsm_0 == 1) && (_source_stream_conv2d_24_source_7_pat_count_0 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_7_pat_cur_offset_1 <= _source_stream_conv2d_24_source_7_pat_cur_offset_1 + _source_stream_conv2d_24_source_7_pat_stride_buf_1;
        _source_stream_conv2d_24_source_7_pat_count_1 <= _source_stream_conv2d_24_source_7_pat_count_1 - 1;
      end 
      if((_stream_conv2d_24_source_7_source_pat_fsm_0 == 1) && (_source_stream_conv2d_24_source_7_pat_count_0 == 0) && (_source_stream_conv2d_24_source_7_pat_count_1 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_7_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_24_source_7_pat_count_1 <= _source_stream_conv2d_24_source_7_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_24_source_7_source_pat_fsm_0 == 1) && ((_source_stream_conv2d_24_source_7_pat_count_0 == 0) && (_source_stream_conv2d_24_source_7_pat_count_1 == 0)) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_7_pat_cur_offset_2 <= _source_stream_conv2d_24_source_7_pat_cur_offset_2 + _source_stream_conv2d_24_source_7_pat_stride_buf_2;
        _source_stream_conv2d_24_source_7_pat_count_2 <= _source_stream_conv2d_24_source_7_pat_count_2 - 1;
      end 
      if((_stream_conv2d_24_source_7_source_pat_fsm_0 == 1) && ((_source_stream_conv2d_24_source_7_pat_count_0 == 0) && (_source_stream_conv2d_24_source_7_pat_count_1 == 0)) && (_source_stream_conv2d_24_source_7_pat_count_2 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_7_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_24_source_7_pat_count_2 <= _source_stream_conv2d_24_source_7_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_24_source_7_source_pat_fsm_0 == 1) && ((_source_stream_conv2d_24_source_7_pat_count_0 == 0) && (_source_stream_conv2d_24_source_7_pat_count_1 == 0) && (_source_stream_conv2d_24_source_7_pat_count_2 == 0)) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_7_pat_cur_offset_3 <= _source_stream_conv2d_24_source_7_pat_cur_offset_3 + _source_stream_conv2d_24_source_7_pat_stride_buf_3;
        _source_stream_conv2d_24_source_7_pat_count_3 <= _source_stream_conv2d_24_source_7_pat_count_3 - 1;
      end 
      if((_stream_conv2d_24_source_7_source_pat_fsm_0 == 1) && ((_source_stream_conv2d_24_source_7_pat_count_0 == 0) && (_source_stream_conv2d_24_source_7_pat_count_1 == 0) && (_source_stream_conv2d_24_source_7_pat_count_2 == 0)) && (_source_stream_conv2d_24_source_7_pat_count_3 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_7_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_24_source_7_pat_count_3 <= _source_stream_conv2d_24_source_7_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_24_source_7_source_pat_fsm_0 == 1) && _stream_conv2d_24_source_stop && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_7_source_ram_renable <= 0;
        _stream_conv2d_24_source_7_idle <= 1;
      end 
      if((_stream_conv2d_24_source_7_source_pat_fsm_0 == 2) && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_7_source_ram_renable <= 0;
        _stream_conv2d_24_source_7_idle <= 1;
      end 
      if(_set_flag_406) begin
        _stream_conv2d_24_parameter_8_next_parameter_data <= cparam_conv2d_24_scale_scala;
      end 
      if(_stream_conv2d_24_source_start) begin
        __variable_wdata_326 <= _stream_conv2d_24_parameter_8_next_parameter_data;
      end 
      if(_set_flag_407) begin
        _stream_conv2d_24_source_9_source_mode <= 5'b10;
        _stream_conv2d_24_source_9_source_offset <= (cparam_conv2d_24_scale_num == 1)? 0 : conv2d_24_och_count_buf;
      end 
      if(_set_flag_407) begin
        _source_stream_conv2d_24_source_9_pat_size_0 <= cparam_conv2d_24_stream_reduce_size;
        _source_stream_conv2d_24_source_9_pat_stride_0 <= 0;
      end 
      if(_set_flag_407) begin
        _source_stream_conv2d_24_source_9_pat_size_1 <= conv2d_24_next_stream_num_ops;
        _source_stream_conv2d_24_source_9_pat_stride_1 <= (cparam_conv2d_24_scale_num == 1)? 0 : 1;
      end 
      if(_set_flag_407) begin
        _source_stream_conv2d_24_source_9_pat_size_2 <= 1;
        _source_stream_conv2d_24_source_9_pat_stride_2 <= 0;
      end 
      if(_set_flag_407) begin
        _source_stream_conv2d_24_source_9_pat_size_3 <= 1;
        _source_stream_conv2d_24_source_9_pat_stride_3 <= 0;
      end 
      if(_set_flag_407) begin
        _stream_conv2d_24_source_9_source_sel <= 2;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_9_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_9_source_offset_buf <= _stream_conv2d_24_source_9_source_offset;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_9_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_9_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_9_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_9_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_9_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_9_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_9_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_9_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_9_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_9_pat_count_0 <= _source_stream_conv2d_24_source_9_pat_size_0 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_9_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_9_pat_count_1 <= _source_stream_conv2d_24_source_9_pat_size_1 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_9_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_9_pat_count_2 <= _source_stream_conv2d_24_source_9_pat_size_2 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_9_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_9_pat_count_3 <= _source_stream_conv2d_24_source_9_pat_size_3 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_9_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_9_pat_size_buf_0 <= _source_stream_conv2d_24_source_9_pat_size_0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_9_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_9_pat_size_buf_1 <= _source_stream_conv2d_24_source_9_pat_size_1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_9_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_9_pat_size_buf_2 <= _source_stream_conv2d_24_source_9_pat_size_2;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_9_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_9_pat_size_buf_3 <= _source_stream_conv2d_24_source_9_pat_size_3;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_9_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_9_pat_stride_buf_0 <= _source_stream_conv2d_24_source_9_pat_stride_0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_9_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_9_pat_stride_buf_1 <= _source_stream_conv2d_24_source_9_pat_stride_1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_9_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_9_pat_stride_buf_2 <= _source_stream_conv2d_24_source_9_pat_stride_2;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_9_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_9_pat_stride_buf_3 <= _source_stream_conv2d_24_source_9_pat_stride_3;
      end 
      if(_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_busy && _stream_conv2d_24_is_root) begin
        __variable_wdata_327 <= _stream_conv2d_24_source_9_source_ram_rdata;
      end 
      if((_stream_conv2d_24_source_9_source_pat_fsm_1 == 1) && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_9_idle <= 0;
        _stream_conv2d_24_source_9_source_ram_raddr <= _stream_conv2d_24_source_9_source_pat_all_offset;
        _stream_conv2d_24_source_9_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_24_source_9_source_pat_fsm_1 == 1) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_9_pat_cur_offset_0 <= _source_stream_conv2d_24_source_9_pat_cur_offset_0 + _source_stream_conv2d_24_source_9_pat_stride_buf_0;
        _source_stream_conv2d_24_source_9_pat_count_0 <= _source_stream_conv2d_24_source_9_pat_count_0 - 1;
      end 
      if((_stream_conv2d_24_source_9_source_pat_fsm_1 == 1) && (_source_stream_conv2d_24_source_9_pat_count_0 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_9_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_24_source_9_pat_count_0 <= _source_stream_conv2d_24_source_9_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_24_source_9_source_pat_fsm_1 == 1) && (_source_stream_conv2d_24_source_9_pat_count_0 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_9_pat_cur_offset_1 <= _source_stream_conv2d_24_source_9_pat_cur_offset_1 + _source_stream_conv2d_24_source_9_pat_stride_buf_1;
        _source_stream_conv2d_24_source_9_pat_count_1 <= _source_stream_conv2d_24_source_9_pat_count_1 - 1;
      end 
      if((_stream_conv2d_24_source_9_source_pat_fsm_1 == 1) && (_source_stream_conv2d_24_source_9_pat_count_0 == 0) && (_source_stream_conv2d_24_source_9_pat_count_1 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_9_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_24_source_9_pat_count_1 <= _source_stream_conv2d_24_source_9_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_24_source_9_source_pat_fsm_1 == 1) && ((_source_stream_conv2d_24_source_9_pat_count_0 == 0) && (_source_stream_conv2d_24_source_9_pat_count_1 == 0)) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_9_pat_cur_offset_2 <= _source_stream_conv2d_24_source_9_pat_cur_offset_2 + _source_stream_conv2d_24_source_9_pat_stride_buf_2;
        _source_stream_conv2d_24_source_9_pat_count_2 <= _source_stream_conv2d_24_source_9_pat_count_2 - 1;
      end 
      if((_stream_conv2d_24_source_9_source_pat_fsm_1 == 1) && ((_source_stream_conv2d_24_source_9_pat_count_0 == 0) && (_source_stream_conv2d_24_source_9_pat_count_1 == 0)) && (_source_stream_conv2d_24_source_9_pat_count_2 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_9_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_24_source_9_pat_count_2 <= _source_stream_conv2d_24_source_9_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_24_source_9_source_pat_fsm_1 == 1) && ((_source_stream_conv2d_24_source_9_pat_count_0 == 0) && (_source_stream_conv2d_24_source_9_pat_count_1 == 0) && (_source_stream_conv2d_24_source_9_pat_count_2 == 0)) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_9_pat_cur_offset_3 <= _source_stream_conv2d_24_source_9_pat_cur_offset_3 + _source_stream_conv2d_24_source_9_pat_stride_buf_3;
        _source_stream_conv2d_24_source_9_pat_count_3 <= _source_stream_conv2d_24_source_9_pat_count_3 - 1;
      end 
      if((_stream_conv2d_24_source_9_source_pat_fsm_1 == 1) && ((_source_stream_conv2d_24_source_9_pat_count_0 == 0) && (_source_stream_conv2d_24_source_9_pat_count_1 == 0) && (_source_stream_conv2d_24_source_9_pat_count_2 == 0)) && (_source_stream_conv2d_24_source_9_pat_count_3 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_9_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_24_source_9_pat_count_3 <= _source_stream_conv2d_24_source_9_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_24_source_9_source_pat_fsm_1 == 1) && _stream_conv2d_24_source_stop && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_9_source_ram_renable <= 0;
        _stream_conv2d_24_source_9_idle <= 1;
      end 
      if((_stream_conv2d_24_source_9_source_pat_fsm_1 == 2) && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_9_source_ram_renable <= 0;
        _stream_conv2d_24_source_9_idle <= 1;
      end 
      if(_set_flag_420) begin
        _stream_conv2d_24_parameter_10_next_parameter_data <= 1;
      end 
      if(_stream_conv2d_24_source_start) begin
        __variable_wdata_333 <= _stream_conv2d_24_parameter_10_next_parameter_data;
      end 
      if(_set_flag_421) begin
        _stream_conv2d_24_source_11_source_mode <= 5'b0;
        _stream_conv2d_24_source_11_source_empty_data <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_stream_oready && !(|(_stream_conv2d_24_source_11_source_mode & 5'b0))) begin
        _stream_conv2d_24_source_11_idle <= 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_stream_oready && !(|(_stream_conv2d_24_source_11_source_mode & 5'b0)) && _stream_conv2d_24_is_root) begin
        __variable_wdata_334 <= _stream_conv2d_24_source_11_source_empty_data;
      end 
      if(_set_flag_422) begin
        _stream_conv2d_24_parameter_12_next_parameter_data <= 1;
      end 
      if(_stream_conv2d_24_source_start) begin
        __variable_wdata_340 <= _stream_conv2d_24_parameter_12_next_parameter_data;
      end 
      if(_set_flag_423) begin
        _stream_conv2d_24_source_13_source_mode <= 5'b0;
        _stream_conv2d_24_source_13_source_empty_data <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_stream_oready && !(|(_stream_conv2d_24_source_13_source_mode & 5'b0))) begin
        _stream_conv2d_24_source_13_idle <= 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_stream_oready && !(|(_stream_conv2d_24_source_13_source_mode & 5'b0)) && _stream_conv2d_24_is_root) begin
        __variable_wdata_341 <= _stream_conv2d_24_source_13_source_empty_data;
      end 
      if(_set_flag_424) begin
        _stream_conv2d_24_parameter_14_next_parameter_data <= 1;
      end 
      if(_stream_conv2d_24_source_start) begin
        __variable_wdata_347 <= _stream_conv2d_24_parameter_14_next_parameter_data;
      end 
      if(_set_flag_425) begin
        _stream_conv2d_24_source_15_source_mode <= 5'b0;
        _stream_conv2d_24_source_15_source_empty_data <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_stream_oready && !(|(_stream_conv2d_24_source_15_source_mode & 5'b0))) begin
        _stream_conv2d_24_source_15_idle <= 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_stream_oready && !(|(_stream_conv2d_24_source_15_source_mode & 5'b0)) && _stream_conv2d_24_is_root) begin
        __variable_wdata_348 <= _stream_conv2d_24_source_15_source_empty_data;
      end 
      if(_set_flag_426) begin
        _stream_conv2d_24_parameter_16_next_parameter_data <= cparam_conv2d_24_cshamt_mul_value;
      end 
      if(_stream_conv2d_24_source_start) begin
        __variable_wdata_354 <= _stream_conv2d_24_parameter_16_next_parameter_data;
      end 
      if(_set_flag_427) begin
        _stream_conv2d_24_parameter_17_next_parameter_data <= cparam_conv2d_24_cshamt_sum_value;
      end 
      if(_stream_conv2d_24_source_start) begin
        __variable_wdata_355 <= _stream_conv2d_24_parameter_17_next_parameter_data;
      end 
      if(_set_flag_428) begin
        _stream_conv2d_24_parameter_18_next_parameter_data <= cparam_conv2d_24_cshamt_out_value;
      end 
      if(_stream_conv2d_24_source_start) begin
        __variable_wdata_356 <= _stream_conv2d_24_parameter_18_next_parameter_data;
      end 
      if(_set_flag_429) begin
        _stream_conv2d_24_parameter_19_next_parameter_data <= cparam_conv2d_24_act_func_index;
      end 
      if(_stream_conv2d_24_source_start) begin
        __variable_wdata_357 <= _stream_conv2d_24_parameter_19_next_parameter_data;
      end 
      if(_set_flag_430) begin
        _stream_conv2d_24_source_20_source_mode <= 5'b10;
        _stream_conv2d_24_source_20_source_offset <= conv2d_24_stream_act_local_0 + conv2d_24_act_page_comp_offset_buf_0;
      end 
      if(_set_flag_430) begin
        _source_stream_conv2d_24_source_20_pat_size_0 <= cparam_conv2d_24_stream_reduce_size;
        _source_stream_conv2d_24_source_20_pat_stride_0 <= 1;
      end 
      if(_set_flag_430) begin
        _source_stream_conv2d_24_source_20_pat_size_1 <= conv2d_24_next_stream_num_ops;
        _source_stream_conv2d_24_source_20_pat_stride_1 <= 0;
      end 
      if(_set_flag_430) begin
        _source_stream_conv2d_24_source_20_pat_size_2 <= 1;
        _source_stream_conv2d_24_source_20_pat_stride_2 <= 0;
      end 
      if(_set_flag_430) begin
        _source_stream_conv2d_24_source_20_pat_size_3 <= 1;
        _source_stream_conv2d_24_source_20_pat_stride_3 <= 0;
      end 
      if(_set_flag_430) begin
        _stream_conv2d_24_source_20_source_sel <= 3;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_20_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_20_source_offset_buf <= _stream_conv2d_24_source_20_source_offset;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_20_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_20_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_20_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_20_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_20_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_20_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_20_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_20_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_20_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_20_pat_count_0 <= _source_stream_conv2d_24_source_20_pat_size_0 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_20_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_20_pat_count_1 <= _source_stream_conv2d_24_source_20_pat_size_1 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_20_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_20_pat_count_2 <= _source_stream_conv2d_24_source_20_pat_size_2 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_20_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_20_pat_count_3 <= _source_stream_conv2d_24_source_20_pat_size_3 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_20_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_20_pat_size_buf_0 <= _source_stream_conv2d_24_source_20_pat_size_0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_20_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_20_pat_size_buf_1 <= _source_stream_conv2d_24_source_20_pat_size_1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_20_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_20_pat_size_buf_2 <= _source_stream_conv2d_24_source_20_pat_size_2;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_20_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_20_pat_size_buf_3 <= _source_stream_conv2d_24_source_20_pat_size_3;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_20_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_20_pat_stride_buf_0 <= _source_stream_conv2d_24_source_20_pat_stride_0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_20_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_20_pat_stride_buf_1 <= _source_stream_conv2d_24_source_20_pat_stride_1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_20_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_20_pat_stride_buf_2 <= _source_stream_conv2d_24_source_20_pat_stride_2;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_20_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_20_pat_stride_buf_3 <= _source_stream_conv2d_24_source_20_pat_stride_3;
      end 
      if(_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_busy && _stream_conv2d_24_is_root) begin
        __variable_wdata_358 <= _stream_conv2d_24_source_20_source_ram_rdata;
      end 
      if((_stream_conv2d_24_source_20_source_pat_fsm_2 == 1) && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_20_idle <= 0;
        _stream_conv2d_24_source_20_source_ram_raddr <= _stream_conv2d_24_source_20_source_pat_all_offset;
        _stream_conv2d_24_source_20_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_24_source_20_source_pat_fsm_2 == 1) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_20_pat_cur_offset_0 <= _source_stream_conv2d_24_source_20_pat_cur_offset_0 + _source_stream_conv2d_24_source_20_pat_stride_buf_0;
        _source_stream_conv2d_24_source_20_pat_count_0 <= _source_stream_conv2d_24_source_20_pat_count_0 - 1;
      end 
      if((_stream_conv2d_24_source_20_source_pat_fsm_2 == 1) && (_source_stream_conv2d_24_source_20_pat_count_0 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_20_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_24_source_20_pat_count_0 <= _source_stream_conv2d_24_source_20_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_24_source_20_source_pat_fsm_2 == 1) && (_source_stream_conv2d_24_source_20_pat_count_0 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_20_pat_cur_offset_1 <= _source_stream_conv2d_24_source_20_pat_cur_offset_1 + _source_stream_conv2d_24_source_20_pat_stride_buf_1;
        _source_stream_conv2d_24_source_20_pat_count_1 <= _source_stream_conv2d_24_source_20_pat_count_1 - 1;
      end 
      if((_stream_conv2d_24_source_20_source_pat_fsm_2 == 1) && (_source_stream_conv2d_24_source_20_pat_count_0 == 0) && (_source_stream_conv2d_24_source_20_pat_count_1 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_20_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_24_source_20_pat_count_1 <= _source_stream_conv2d_24_source_20_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_24_source_20_source_pat_fsm_2 == 1) && ((_source_stream_conv2d_24_source_20_pat_count_0 == 0) && (_source_stream_conv2d_24_source_20_pat_count_1 == 0)) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_20_pat_cur_offset_2 <= _source_stream_conv2d_24_source_20_pat_cur_offset_2 + _source_stream_conv2d_24_source_20_pat_stride_buf_2;
        _source_stream_conv2d_24_source_20_pat_count_2 <= _source_stream_conv2d_24_source_20_pat_count_2 - 1;
      end 
      if((_stream_conv2d_24_source_20_source_pat_fsm_2 == 1) && ((_source_stream_conv2d_24_source_20_pat_count_0 == 0) && (_source_stream_conv2d_24_source_20_pat_count_1 == 0)) && (_source_stream_conv2d_24_source_20_pat_count_2 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_20_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_24_source_20_pat_count_2 <= _source_stream_conv2d_24_source_20_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_24_source_20_source_pat_fsm_2 == 1) && ((_source_stream_conv2d_24_source_20_pat_count_0 == 0) && (_source_stream_conv2d_24_source_20_pat_count_1 == 0) && (_source_stream_conv2d_24_source_20_pat_count_2 == 0)) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_20_pat_cur_offset_3 <= _source_stream_conv2d_24_source_20_pat_cur_offset_3 + _source_stream_conv2d_24_source_20_pat_stride_buf_3;
        _source_stream_conv2d_24_source_20_pat_count_3 <= _source_stream_conv2d_24_source_20_pat_count_3 - 1;
      end 
      if((_stream_conv2d_24_source_20_source_pat_fsm_2 == 1) && ((_source_stream_conv2d_24_source_20_pat_count_0 == 0) && (_source_stream_conv2d_24_source_20_pat_count_1 == 0) && (_source_stream_conv2d_24_source_20_pat_count_2 == 0)) && (_source_stream_conv2d_24_source_20_pat_count_3 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_20_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_24_source_20_pat_count_3 <= _source_stream_conv2d_24_source_20_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_24_source_20_source_pat_fsm_2 == 1) && _stream_conv2d_24_source_stop && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_20_source_ram_renable <= 0;
        _stream_conv2d_24_source_20_idle <= 1;
      end 
      if((_stream_conv2d_24_source_20_source_pat_fsm_2 == 2) && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_20_source_ram_renable <= 0;
        _stream_conv2d_24_source_20_idle <= 1;
      end 
      if(_set_flag_443) begin
        _stream_conv2d_24_source_21_source_mode <= 5'b10;
        _stream_conv2d_24_source_21_source_offset <= conv2d_24_stream_act_local_1 + conv2d_24_act_page_comp_offset_buf_0;
      end 
      if(_set_flag_443) begin
        _source_stream_conv2d_24_source_21_pat_size_0 <= cparam_conv2d_24_stream_reduce_size;
        _source_stream_conv2d_24_source_21_pat_stride_0 <= 1;
      end 
      if(_set_flag_443) begin
        _source_stream_conv2d_24_source_21_pat_size_1 <= conv2d_24_next_stream_num_ops;
        _source_stream_conv2d_24_source_21_pat_stride_1 <= 0;
      end 
      if(_set_flag_443) begin
        _source_stream_conv2d_24_source_21_pat_size_2 <= 1;
        _source_stream_conv2d_24_source_21_pat_stride_2 <= 0;
      end 
      if(_set_flag_443) begin
        _source_stream_conv2d_24_source_21_pat_size_3 <= 1;
        _source_stream_conv2d_24_source_21_pat_stride_3 <= 0;
      end 
      if(_set_flag_443) begin
        _stream_conv2d_24_source_21_source_sel <= 4;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_21_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_21_source_offset_buf <= _stream_conv2d_24_source_21_source_offset;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_21_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_21_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_21_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_21_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_21_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_21_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_21_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_21_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_21_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_21_pat_count_0 <= _source_stream_conv2d_24_source_21_pat_size_0 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_21_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_21_pat_count_1 <= _source_stream_conv2d_24_source_21_pat_size_1 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_21_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_21_pat_count_2 <= _source_stream_conv2d_24_source_21_pat_size_2 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_21_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_21_pat_count_3 <= _source_stream_conv2d_24_source_21_pat_size_3 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_21_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_21_pat_size_buf_0 <= _source_stream_conv2d_24_source_21_pat_size_0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_21_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_21_pat_size_buf_1 <= _source_stream_conv2d_24_source_21_pat_size_1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_21_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_21_pat_size_buf_2 <= _source_stream_conv2d_24_source_21_pat_size_2;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_21_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_21_pat_size_buf_3 <= _source_stream_conv2d_24_source_21_pat_size_3;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_21_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_21_pat_stride_buf_0 <= _source_stream_conv2d_24_source_21_pat_stride_0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_21_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_21_pat_stride_buf_1 <= _source_stream_conv2d_24_source_21_pat_stride_1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_21_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_21_pat_stride_buf_2 <= _source_stream_conv2d_24_source_21_pat_stride_2;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_21_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_21_pat_stride_buf_3 <= _source_stream_conv2d_24_source_21_pat_stride_3;
      end 
      if(_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_busy && _stream_conv2d_24_is_root) begin
        __variable_wdata_359 <= _stream_conv2d_24_source_21_source_ram_rdata;
      end 
      if((_stream_conv2d_24_source_21_source_pat_fsm_3 == 1) && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_21_idle <= 0;
        _stream_conv2d_24_source_21_source_ram_raddr <= _stream_conv2d_24_source_21_source_pat_all_offset;
        _stream_conv2d_24_source_21_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_24_source_21_source_pat_fsm_3 == 1) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_21_pat_cur_offset_0 <= _source_stream_conv2d_24_source_21_pat_cur_offset_0 + _source_stream_conv2d_24_source_21_pat_stride_buf_0;
        _source_stream_conv2d_24_source_21_pat_count_0 <= _source_stream_conv2d_24_source_21_pat_count_0 - 1;
      end 
      if((_stream_conv2d_24_source_21_source_pat_fsm_3 == 1) && (_source_stream_conv2d_24_source_21_pat_count_0 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_21_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_24_source_21_pat_count_0 <= _source_stream_conv2d_24_source_21_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_24_source_21_source_pat_fsm_3 == 1) && (_source_stream_conv2d_24_source_21_pat_count_0 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_21_pat_cur_offset_1 <= _source_stream_conv2d_24_source_21_pat_cur_offset_1 + _source_stream_conv2d_24_source_21_pat_stride_buf_1;
        _source_stream_conv2d_24_source_21_pat_count_1 <= _source_stream_conv2d_24_source_21_pat_count_1 - 1;
      end 
      if((_stream_conv2d_24_source_21_source_pat_fsm_3 == 1) && (_source_stream_conv2d_24_source_21_pat_count_0 == 0) && (_source_stream_conv2d_24_source_21_pat_count_1 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_21_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_24_source_21_pat_count_1 <= _source_stream_conv2d_24_source_21_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_24_source_21_source_pat_fsm_3 == 1) && ((_source_stream_conv2d_24_source_21_pat_count_0 == 0) && (_source_stream_conv2d_24_source_21_pat_count_1 == 0)) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_21_pat_cur_offset_2 <= _source_stream_conv2d_24_source_21_pat_cur_offset_2 + _source_stream_conv2d_24_source_21_pat_stride_buf_2;
        _source_stream_conv2d_24_source_21_pat_count_2 <= _source_stream_conv2d_24_source_21_pat_count_2 - 1;
      end 
      if((_stream_conv2d_24_source_21_source_pat_fsm_3 == 1) && ((_source_stream_conv2d_24_source_21_pat_count_0 == 0) && (_source_stream_conv2d_24_source_21_pat_count_1 == 0)) && (_source_stream_conv2d_24_source_21_pat_count_2 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_21_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_24_source_21_pat_count_2 <= _source_stream_conv2d_24_source_21_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_24_source_21_source_pat_fsm_3 == 1) && ((_source_stream_conv2d_24_source_21_pat_count_0 == 0) && (_source_stream_conv2d_24_source_21_pat_count_1 == 0) && (_source_stream_conv2d_24_source_21_pat_count_2 == 0)) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_21_pat_cur_offset_3 <= _source_stream_conv2d_24_source_21_pat_cur_offset_3 + _source_stream_conv2d_24_source_21_pat_stride_buf_3;
        _source_stream_conv2d_24_source_21_pat_count_3 <= _source_stream_conv2d_24_source_21_pat_count_3 - 1;
      end 
      if((_stream_conv2d_24_source_21_source_pat_fsm_3 == 1) && ((_source_stream_conv2d_24_source_21_pat_count_0 == 0) && (_source_stream_conv2d_24_source_21_pat_count_1 == 0) && (_source_stream_conv2d_24_source_21_pat_count_2 == 0)) && (_source_stream_conv2d_24_source_21_pat_count_3 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_21_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_24_source_21_pat_count_3 <= _source_stream_conv2d_24_source_21_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_24_source_21_source_pat_fsm_3 == 1) && _stream_conv2d_24_source_stop && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_21_source_ram_renable <= 0;
        _stream_conv2d_24_source_21_idle <= 1;
      end 
      if((_stream_conv2d_24_source_21_source_pat_fsm_3 == 2) && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_21_source_ram_renable <= 0;
        _stream_conv2d_24_source_21_idle <= 1;
      end 
      if(_set_flag_456) begin
        _stream_conv2d_24_source_22_source_mode <= 5'b10;
        _stream_conv2d_24_source_22_source_offset <= conv2d_24_stream_act_local_2 + conv2d_24_act_page_comp_offset_buf_0;
      end 
      if(_set_flag_456) begin
        _source_stream_conv2d_24_source_22_pat_size_0 <= cparam_conv2d_24_stream_reduce_size;
        _source_stream_conv2d_24_source_22_pat_stride_0 <= 1;
      end 
      if(_set_flag_456) begin
        _source_stream_conv2d_24_source_22_pat_size_1 <= conv2d_24_next_stream_num_ops;
        _source_stream_conv2d_24_source_22_pat_stride_1 <= 0;
      end 
      if(_set_flag_456) begin
        _source_stream_conv2d_24_source_22_pat_size_2 <= 1;
        _source_stream_conv2d_24_source_22_pat_stride_2 <= 0;
      end 
      if(_set_flag_456) begin
        _source_stream_conv2d_24_source_22_pat_size_3 <= 1;
        _source_stream_conv2d_24_source_22_pat_stride_3 <= 0;
      end 
      if(_set_flag_456) begin
        _stream_conv2d_24_source_22_source_sel <= 5;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_22_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_22_source_offset_buf <= _stream_conv2d_24_source_22_source_offset;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_22_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_22_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_22_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_22_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_22_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_22_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_22_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_22_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_22_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_22_pat_count_0 <= _source_stream_conv2d_24_source_22_pat_size_0 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_22_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_22_pat_count_1 <= _source_stream_conv2d_24_source_22_pat_size_1 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_22_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_22_pat_count_2 <= _source_stream_conv2d_24_source_22_pat_size_2 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_22_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_22_pat_count_3 <= _source_stream_conv2d_24_source_22_pat_size_3 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_22_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_22_pat_size_buf_0 <= _source_stream_conv2d_24_source_22_pat_size_0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_22_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_22_pat_size_buf_1 <= _source_stream_conv2d_24_source_22_pat_size_1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_22_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_22_pat_size_buf_2 <= _source_stream_conv2d_24_source_22_pat_size_2;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_22_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_22_pat_size_buf_3 <= _source_stream_conv2d_24_source_22_pat_size_3;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_22_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_22_pat_stride_buf_0 <= _source_stream_conv2d_24_source_22_pat_stride_0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_22_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_22_pat_stride_buf_1 <= _source_stream_conv2d_24_source_22_pat_stride_1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_22_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_22_pat_stride_buf_2 <= _source_stream_conv2d_24_source_22_pat_stride_2;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_22_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_22_pat_stride_buf_3 <= _source_stream_conv2d_24_source_22_pat_stride_3;
      end 
      if(_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_busy && _stream_conv2d_24_is_root) begin
        __variable_wdata_360 <= _stream_conv2d_24_source_22_source_ram_rdata;
      end 
      if((_stream_conv2d_24_source_22_source_pat_fsm_4 == 1) && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_22_idle <= 0;
        _stream_conv2d_24_source_22_source_ram_raddr <= _stream_conv2d_24_source_22_source_pat_all_offset;
        _stream_conv2d_24_source_22_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_24_source_22_source_pat_fsm_4 == 1) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_22_pat_cur_offset_0 <= _source_stream_conv2d_24_source_22_pat_cur_offset_0 + _source_stream_conv2d_24_source_22_pat_stride_buf_0;
        _source_stream_conv2d_24_source_22_pat_count_0 <= _source_stream_conv2d_24_source_22_pat_count_0 - 1;
      end 
      if((_stream_conv2d_24_source_22_source_pat_fsm_4 == 1) && (_source_stream_conv2d_24_source_22_pat_count_0 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_22_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_24_source_22_pat_count_0 <= _source_stream_conv2d_24_source_22_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_24_source_22_source_pat_fsm_4 == 1) && (_source_stream_conv2d_24_source_22_pat_count_0 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_22_pat_cur_offset_1 <= _source_stream_conv2d_24_source_22_pat_cur_offset_1 + _source_stream_conv2d_24_source_22_pat_stride_buf_1;
        _source_stream_conv2d_24_source_22_pat_count_1 <= _source_stream_conv2d_24_source_22_pat_count_1 - 1;
      end 
      if((_stream_conv2d_24_source_22_source_pat_fsm_4 == 1) && (_source_stream_conv2d_24_source_22_pat_count_0 == 0) && (_source_stream_conv2d_24_source_22_pat_count_1 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_22_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_24_source_22_pat_count_1 <= _source_stream_conv2d_24_source_22_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_24_source_22_source_pat_fsm_4 == 1) && ((_source_stream_conv2d_24_source_22_pat_count_0 == 0) && (_source_stream_conv2d_24_source_22_pat_count_1 == 0)) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_22_pat_cur_offset_2 <= _source_stream_conv2d_24_source_22_pat_cur_offset_2 + _source_stream_conv2d_24_source_22_pat_stride_buf_2;
        _source_stream_conv2d_24_source_22_pat_count_2 <= _source_stream_conv2d_24_source_22_pat_count_2 - 1;
      end 
      if((_stream_conv2d_24_source_22_source_pat_fsm_4 == 1) && ((_source_stream_conv2d_24_source_22_pat_count_0 == 0) && (_source_stream_conv2d_24_source_22_pat_count_1 == 0)) && (_source_stream_conv2d_24_source_22_pat_count_2 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_22_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_24_source_22_pat_count_2 <= _source_stream_conv2d_24_source_22_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_24_source_22_source_pat_fsm_4 == 1) && ((_source_stream_conv2d_24_source_22_pat_count_0 == 0) && (_source_stream_conv2d_24_source_22_pat_count_1 == 0) && (_source_stream_conv2d_24_source_22_pat_count_2 == 0)) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_22_pat_cur_offset_3 <= _source_stream_conv2d_24_source_22_pat_cur_offset_3 + _source_stream_conv2d_24_source_22_pat_stride_buf_3;
        _source_stream_conv2d_24_source_22_pat_count_3 <= _source_stream_conv2d_24_source_22_pat_count_3 - 1;
      end 
      if((_stream_conv2d_24_source_22_source_pat_fsm_4 == 1) && ((_source_stream_conv2d_24_source_22_pat_count_0 == 0) && (_source_stream_conv2d_24_source_22_pat_count_1 == 0) && (_source_stream_conv2d_24_source_22_pat_count_2 == 0)) && (_source_stream_conv2d_24_source_22_pat_count_3 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_22_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_24_source_22_pat_count_3 <= _source_stream_conv2d_24_source_22_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_24_source_22_source_pat_fsm_4 == 1) && _stream_conv2d_24_source_stop && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_22_source_ram_renable <= 0;
        _stream_conv2d_24_source_22_idle <= 1;
      end 
      if((_stream_conv2d_24_source_22_source_pat_fsm_4 == 2) && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_22_source_ram_renable <= 0;
        _stream_conv2d_24_source_22_idle <= 1;
      end 
      if(_set_flag_469) begin
        _stream_conv2d_24_source_23_source_mode <= 5'b10;
        _stream_conv2d_24_source_23_source_offset <= conv2d_24_stream_act_local_3 + conv2d_24_act_page_comp_offset_buf_1;
      end 
      if(_set_flag_469) begin
        _source_stream_conv2d_24_source_23_pat_size_0 <= cparam_conv2d_24_stream_reduce_size;
        _source_stream_conv2d_24_source_23_pat_stride_0 <= 1;
      end 
      if(_set_flag_469) begin
        _source_stream_conv2d_24_source_23_pat_size_1 <= conv2d_24_next_stream_num_ops;
        _source_stream_conv2d_24_source_23_pat_stride_1 <= 0;
      end 
      if(_set_flag_469) begin
        _source_stream_conv2d_24_source_23_pat_size_2 <= 1;
        _source_stream_conv2d_24_source_23_pat_stride_2 <= 0;
      end 
      if(_set_flag_469) begin
        _source_stream_conv2d_24_source_23_pat_size_3 <= 1;
        _source_stream_conv2d_24_source_23_pat_stride_3 <= 0;
      end 
      if(_set_flag_469) begin
        _stream_conv2d_24_source_23_source_sel <= 6;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_23_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_23_source_offset_buf <= _stream_conv2d_24_source_23_source_offset;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_23_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_23_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_23_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_23_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_23_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_23_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_23_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_23_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_23_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_23_pat_count_0 <= _source_stream_conv2d_24_source_23_pat_size_0 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_23_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_23_pat_count_1 <= _source_stream_conv2d_24_source_23_pat_size_1 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_23_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_23_pat_count_2 <= _source_stream_conv2d_24_source_23_pat_size_2 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_23_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_23_pat_count_3 <= _source_stream_conv2d_24_source_23_pat_size_3 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_23_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_23_pat_size_buf_0 <= _source_stream_conv2d_24_source_23_pat_size_0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_23_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_23_pat_size_buf_1 <= _source_stream_conv2d_24_source_23_pat_size_1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_23_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_23_pat_size_buf_2 <= _source_stream_conv2d_24_source_23_pat_size_2;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_23_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_23_pat_size_buf_3 <= _source_stream_conv2d_24_source_23_pat_size_3;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_23_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_23_pat_stride_buf_0 <= _source_stream_conv2d_24_source_23_pat_stride_0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_23_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_23_pat_stride_buf_1 <= _source_stream_conv2d_24_source_23_pat_stride_1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_23_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_23_pat_stride_buf_2 <= _source_stream_conv2d_24_source_23_pat_stride_2;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_23_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_23_pat_stride_buf_3 <= _source_stream_conv2d_24_source_23_pat_stride_3;
      end 
      if(_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_busy && _stream_conv2d_24_is_root) begin
        __variable_wdata_361 <= _stream_conv2d_24_source_23_source_ram_rdata;
      end 
      if((_stream_conv2d_24_source_23_source_pat_fsm_5 == 1) && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_23_idle <= 0;
        _stream_conv2d_24_source_23_source_ram_raddr <= _stream_conv2d_24_source_23_source_pat_all_offset;
        _stream_conv2d_24_source_23_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_24_source_23_source_pat_fsm_5 == 1) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_23_pat_cur_offset_0 <= _source_stream_conv2d_24_source_23_pat_cur_offset_0 + _source_stream_conv2d_24_source_23_pat_stride_buf_0;
        _source_stream_conv2d_24_source_23_pat_count_0 <= _source_stream_conv2d_24_source_23_pat_count_0 - 1;
      end 
      if((_stream_conv2d_24_source_23_source_pat_fsm_5 == 1) && (_source_stream_conv2d_24_source_23_pat_count_0 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_23_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_24_source_23_pat_count_0 <= _source_stream_conv2d_24_source_23_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_24_source_23_source_pat_fsm_5 == 1) && (_source_stream_conv2d_24_source_23_pat_count_0 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_23_pat_cur_offset_1 <= _source_stream_conv2d_24_source_23_pat_cur_offset_1 + _source_stream_conv2d_24_source_23_pat_stride_buf_1;
        _source_stream_conv2d_24_source_23_pat_count_1 <= _source_stream_conv2d_24_source_23_pat_count_1 - 1;
      end 
      if((_stream_conv2d_24_source_23_source_pat_fsm_5 == 1) && (_source_stream_conv2d_24_source_23_pat_count_0 == 0) && (_source_stream_conv2d_24_source_23_pat_count_1 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_23_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_24_source_23_pat_count_1 <= _source_stream_conv2d_24_source_23_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_24_source_23_source_pat_fsm_5 == 1) && ((_source_stream_conv2d_24_source_23_pat_count_0 == 0) && (_source_stream_conv2d_24_source_23_pat_count_1 == 0)) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_23_pat_cur_offset_2 <= _source_stream_conv2d_24_source_23_pat_cur_offset_2 + _source_stream_conv2d_24_source_23_pat_stride_buf_2;
        _source_stream_conv2d_24_source_23_pat_count_2 <= _source_stream_conv2d_24_source_23_pat_count_2 - 1;
      end 
      if((_stream_conv2d_24_source_23_source_pat_fsm_5 == 1) && ((_source_stream_conv2d_24_source_23_pat_count_0 == 0) && (_source_stream_conv2d_24_source_23_pat_count_1 == 0)) && (_source_stream_conv2d_24_source_23_pat_count_2 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_23_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_24_source_23_pat_count_2 <= _source_stream_conv2d_24_source_23_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_24_source_23_source_pat_fsm_5 == 1) && ((_source_stream_conv2d_24_source_23_pat_count_0 == 0) && (_source_stream_conv2d_24_source_23_pat_count_1 == 0) && (_source_stream_conv2d_24_source_23_pat_count_2 == 0)) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_23_pat_cur_offset_3 <= _source_stream_conv2d_24_source_23_pat_cur_offset_3 + _source_stream_conv2d_24_source_23_pat_stride_buf_3;
        _source_stream_conv2d_24_source_23_pat_count_3 <= _source_stream_conv2d_24_source_23_pat_count_3 - 1;
      end 
      if((_stream_conv2d_24_source_23_source_pat_fsm_5 == 1) && ((_source_stream_conv2d_24_source_23_pat_count_0 == 0) && (_source_stream_conv2d_24_source_23_pat_count_1 == 0) && (_source_stream_conv2d_24_source_23_pat_count_2 == 0)) && (_source_stream_conv2d_24_source_23_pat_count_3 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_23_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_24_source_23_pat_count_3 <= _source_stream_conv2d_24_source_23_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_24_source_23_source_pat_fsm_5 == 1) && _stream_conv2d_24_source_stop && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_23_source_ram_renable <= 0;
        _stream_conv2d_24_source_23_idle <= 1;
      end 
      if((_stream_conv2d_24_source_23_source_pat_fsm_5 == 2) && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_23_source_ram_renable <= 0;
        _stream_conv2d_24_source_23_idle <= 1;
      end 
      if(_set_flag_482) begin
        _stream_conv2d_24_source_24_source_mode <= 5'b10;
        _stream_conv2d_24_source_24_source_offset <= conv2d_24_stream_act_local_4 + conv2d_24_act_page_comp_offset_buf_1;
      end 
      if(_set_flag_482) begin
        _source_stream_conv2d_24_source_24_pat_size_0 <= cparam_conv2d_24_stream_reduce_size;
        _source_stream_conv2d_24_source_24_pat_stride_0 <= 1;
      end 
      if(_set_flag_482) begin
        _source_stream_conv2d_24_source_24_pat_size_1 <= conv2d_24_next_stream_num_ops;
        _source_stream_conv2d_24_source_24_pat_stride_1 <= 0;
      end 
      if(_set_flag_482) begin
        _source_stream_conv2d_24_source_24_pat_size_2 <= 1;
        _source_stream_conv2d_24_source_24_pat_stride_2 <= 0;
      end 
      if(_set_flag_482) begin
        _source_stream_conv2d_24_source_24_pat_size_3 <= 1;
        _source_stream_conv2d_24_source_24_pat_stride_3 <= 0;
      end 
      if(_set_flag_482) begin
        _stream_conv2d_24_source_24_source_sel <= 7;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_24_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_24_source_offset_buf <= _stream_conv2d_24_source_24_source_offset;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_24_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_24_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_24_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_24_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_24_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_24_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_24_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_24_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_24_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_24_pat_count_0 <= _source_stream_conv2d_24_source_24_pat_size_0 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_24_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_24_pat_count_1 <= _source_stream_conv2d_24_source_24_pat_size_1 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_24_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_24_pat_count_2 <= _source_stream_conv2d_24_source_24_pat_size_2 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_24_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_24_pat_count_3 <= _source_stream_conv2d_24_source_24_pat_size_3 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_24_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_24_pat_size_buf_0 <= _source_stream_conv2d_24_source_24_pat_size_0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_24_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_24_pat_size_buf_1 <= _source_stream_conv2d_24_source_24_pat_size_1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_24_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_24_pat_size_buf_2 <= _source_stream_conv2d_24_source_24_pat_size_2;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_24_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_24_pat_size_buf_3 <= _source_stream_conv2d_24_source_24_pat_size_3;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_24_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_24_pat_stride_buf_0 <= _source_stream_conv2d_24_source_24_pat_stride_0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_24_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_24_pat_stride_buf_1 <= _source_stream_conv2d_24_source_24_pat_stride_1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_24_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_24_pat_stride_buf_2 <= _source_stream_conv2d_24_source_24_pat_stride_2;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_24_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_24_pat_stride_buf_3 <= _source_stream_conv2d_24_source_24_pat_stride_3;
      end 
      if(_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_busy && _stream_conv2d_24_is_root) begin
        __variable_wdata_362 <= _stream_conv2d_24_source_24_source_ram_rdata;
      end 
      if((_stream_conv2d_24_source_24_source_pat_fsm_6 == 1) && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_24_idle <= 0;
        _stream_conv2d_24_source_24_source_ram_raddr <= _stream_conv2d_24_source_24_source_pat_all_offset;
        _stream_conv2d_24_source_24_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_24_source_24_source_pat_fsm_6 == 1) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_24_pat_cur_offset_0 <= _source_stream_conv2d_24_source_24_pat_cur_offset_0 + _source_stream_conv2d_24_source_24_pat_stride_buf_0;
        _source_stream_conv2d_24_source_24_pat_count_0 <= _source_stream_conv2d_24_source_24_pat_count_0 - 1;
      end 
      if((_stream_conv2d_24_source_24_source_pat_fsm_6 == 1) && (_source_stream_conv2d_24_source_24_pat_count_0 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_24_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_24_source_24_pat_count_0 <= _source_stream_conv2d_24_source_24_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_24_source_24_source_pat_fsm_6 == 1) && (_source_stream_conv2d_24_source_24_pat_count_0 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_24_pat_cur_offset_1 <= _source_stream_conv2d_24_source_24_pat_cur_offset_1 + _source_stream_conv2d_24_source_24_pat_stride_buf_1;
        _source_stream_conv2d_24_source_24_pat_count_1 <= _source_stream_conv2d_24_source_24_pat_count_1 - 1;
      end 
      if((_stream_conv2d_24_source_24_source_pat_fsm_6 == 1) && (_source_stream_conv2d_24_source_24_pat_count_0 == 0) && (_source_stream_conv2d_24_source_24_pat_count_1 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_24_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_24_source_24_pat_count_1 <= _source_stream_conv2d_24_source_24_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_24_source_24_source_pat_fsm_6 == 1) && ((_source_stream_conv2d_24_source_24_pat_count_0 == 0) && (_source_stream_conv2d_24_source_24_pat_count_1 == 0)) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_24_pat_cur_offset_2 <= _source_stream_conv2d_24_source_24_pat_cur_offset_2 + _source_stream_conv2d_24_source_24_pat_stride_buf_2;
        _source_stream_conv2d_24_source_24_pat_count_2 <= _source_stream_conv2d_24_source_24_pat_count_2 - 1;
      end 
      if((_stream_conv2d_24_source_24_source_pat_fsm_6 == 1) && ((_source_stream_conv2d_24_source_24_pat_count_0 == 0) && (_source_stream_conv2d_24_source_24_pat_count_1 == 0)) && (_source_stream_conv2d_24_source_24_pat_count_2 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_24_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_24_source_24_pat_count_2 <= _source_stream_conv2d_24_source_24_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_24_source_24_source_pat_fsm_6 == 1) && ((_source_stream_conv2d_24_source_24_pat_count_0 == 0) && (_source_stream_conv2d_24_source_24_pat_count_1 == 0) && (_source_stream_conv2d_24_source_24_pat_count_2 == 0)) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_24_pat_cur_offset_3 <= _source_stream_conv2d_24_source_24_pat_cur_offset_3 + _source_stream_conv2d_24_source_24_pat_stride_buf_3;
        _source_stream_conv2d_24_source_24_pat_count_3 <= _source_stream_conv2d_24_source_24_pat_count_3 - 1;
      end 
      if((_stream_conv2d_24_source_24_source_pat_fsm_6 == 1) && ((_source_stream_conv2d_24_source_24_pat_count_0 == 0) && (_source_stream_conv2d_24_source_24_pat_count_1 == 0) && (_source_stream_conv2d_24_source_24_pat_count_2 == 0)) && (_source_stream_conv2d_24_source_24_pat_count_3 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_24_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_24_source_24_pat_count_3 <= _source_stream_conv2d_24_source_24_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_24_source_24_source_pat_fsm_6 == 1) && _stream_conv2d_24_source_stop && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_24_source_ram_renable <= 0;
        _stream_conv2d_24_source_24_idle <= 1;
      end 
      if((_stream_conv2d_24_source_24_source_pat_fsm_6 == 2) && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_24_source_ram_renable <= 0;
        _stream_conv2d_24_source_24_idle <= 1;
      end 
      if(_set_flag_495) begin
        _stream_conv2d_24_source_25_source_mode <= 5'b10;
        _stream_conv2d_24_source_25_source_offset <= conv2d_24_stream_act_local_5 + conv2d_24_act_page_comp_offset_buf_1;
      end 
      if(_set_flag_495) begin
        _source_stream_conv2d_24_source_25_pat_size_0 <= cparam_conv2d_24_stream_reduce_size;
        _source_stream_conv2d_24_source_25_pat_stride_0 <= 1;
      end 
      if(_set_flag_495) begin
        _source_stream_conv2d_24_source_25_pat_size_1 <= conv2d_24_next_stream_num_ops;
        _source_stream_conv2d_24_source_25_pat_stride_1 <= 0;
      end 
      if(_set_flag_495) begin
        _source_stream_conv2d_24_source_25_pat_size_2 <= 1;
        _source_stream_conv2d_24_source_25_pat_stride_2 <= 0;
      end 
      if(_set_flag_495) begin
        _source_stream_conv2d_24_source_25_pat_size_3 <= 1;
        _source_stream_conv2d_24_source_25_pat_stride_3 <= 0;
      end 
      if(_set_flag_495) begin
        _stream_conv2d_24_source_25_source_sel <= 8;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_25_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_25_source_offset_buf <= _stream_conv2d_24_source_25_source_offset;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_25_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_25_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_25_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_25_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_25_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_25_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_25_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_25_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_25_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_25_pat_count_0 <= _source_stream_conv2d_24_source_25_pat_size_0 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_25_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_25_pat_count_1 <= _source_stream_conv2d_24_source_25_pat_size_1 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_25_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_25_pat_count_2 <= _source_stream_conv2d_24_source_25_pat_size_2 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_25_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_25_pat_count_3 <= _source_stream_conv2d_24_source_25_pat_size_3 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_25_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_25_pat_size_buf_0 <= _source_stream_conv2d_24_source_25_pat_size_0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_25_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_25_pat_size_buf_1 <= _source_stream_conv2d_24_source_25_pat_size_1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_25_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_25_pat_size_buf_2 <= _source_stream_conv2d_24_source_25_pat_size_2;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_25_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_25_pat_size_buf_3 <= _source_stream_conv2d_24_source_25_pat_size_3;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_25_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_25_pat_stride_buf_0 <= _source_stream_conv2d_24_source_25_pat_stride_0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_25_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_25_pat_stride_buf_1 <= _source_stream_conv2d_24_source_25_pat_stride_1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_25_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_25_pat_stride_buf_2 <= _source_stream_conv2d_24_source_25_pat_stride_2;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_25_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_25_pat_stride_buf_3 <= _source_stream_conv2d_24_source_25_pat_stride_3;
      end 
      if(_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_busy && _stream_conv2d_24_is_root) begin
        __variable_wdata_363 <= _stream_conv2d_24_source_25_source_ram_rdata;
      end 
      if((_stream_conv2d_24_source_25_source_pat_fsm_7 == 1) && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_25_idle <= 0;
        _stream_conv2d_24_source_25_source_ram_raddr <= _stream_conv2d_24_source_25_source_pat_all_offset;
        _stream_conv2d_24_source_25_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_24_source_25_source_pat_fsm_7 == 1) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_25_pat_cur_offset_0 <= _source_stream_conv2d_24_source_25_pat_cur_offset_0 + _source_stream_conv2d_24_source_25_pat_stride_buf_0;
        _source_stream_conv2d_24_source_25_pat_count_0 <= _source_stream_conv2d_24_source_25_pat_count_0 - 1;
      end 
      if((_stream_conv2d_24_source_25_source_pat_fsm_7 == 1) && (_source_stream_conv2d_24_source_25_pat_count_0 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_25_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_24_source_25_pat_count_0 <= _source_stream_conv2d_24_source_25_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_24_source_25_source_pat_fsm_7 == 1) && (_source_stream_conv2d_24_source_25_pat_count_0 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_25_pat_cur_offset_1 <= _source_stream_conv2d_24_source_25_pat_cur_offset_1 + _source_stream_conv2d_24_source_25_pat_stride_buf_1;
        _source_stream_conv2d_24_source_25_pat_count_1 <= _source_stream_conv2d_24_source_25_pat_count_1 - 1;
      end 
      if((_stream_conv2d_24_source_25_source_pat_fsm_7 == 1) && (_source_stream_conv2d_24_source_25_pat_count_0 == 0) && (_source_stream_conv2d_24_source_25_pat_count_1 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_25_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_24_source_25_pat_count_1 <= _source_stream_conv2d_24_source_25_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_24_source_25_source_pat_fsm_7 == 1) && ((_source_stream_conv2d_24_source_25_pat_count_0 == 0) && (_source_stream_conv2d_24_source_25_pat_count_1 == 0)) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_25_pat_cur_offset_2 <= _source_stream_conv2d_24_source_25_pat_cur_offset_2 + _source_stream_conv2d_24_source_25_pat_stride_buf_2;
        _source_stream_conv2d_24_source_25_pat_count_2 <= _source_stream_conv2d_24_source_25_pat_count_2 - 1;
      end 
      if((_stream_conv2d_24_source_25_source_pat_fsm_7 == 1) && ((_source_stream_conv2d_24_source_25_pat_count_0 == 0) && (_source_stream_conv2d_24_source_25_pat_count_1 == 0)) && (_source_stream_conv2d_24_source_25_pat_count_2 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_25_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_24_source_25_pat_count_2 <= _source_stream_conv2d_24_source_25_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_24_source_25_source_pat_fsm_7 == 1) && ((_source_stream_conv2d_24_source_25_pat_count_0 == 0) && (_source_stream_conv2d_24_source_25_pat_count_1 == 0) && (_source_stream_conv2d_24_source_25_pat_count_2 == 0)) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_25_pat_cur_offset_3 <= _source_stream_conv2d_24_source_25_pat_cur_offset_3 + _source_stream_conv2d_24_source_25_pat_stride_buf_3;
        _source_stream_conv2d_24_source_25_pat_count_3 <= _source_stream_conv2d_24_source_25_pat_count_3 - 1;
      end 
      if((_stream_conv2d_24_source_25_source_pat_fsm_7 == 1) && ((_source_stream_conv2d_24_source_25_pat_count_0 == 0) && (_source_stream_conv2d_24_source_25_pat_count_1 == 0) && (_source_stream_conv2d_24_source_25_pat_count_2 == 0)) && (_source_stream_conv2d_24_source_25_pat_count_3 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_25_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_24_source_25_pat_count_3 <= _source_stream_conv2d_24_source_25_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_24_source_25_source_pat_fsm_7 == 1) && _stream_conv2d_24_source_stop && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_25_source_ram_renable <= 0;
        _stream_conv2d_24_source_25_idle <= 1;
      end 
      if((_stream_conv2d_24_source_25_source_pat_fsm_7 == 2) && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_25_source_ram_renable <= 0;
        _stream_conv2d_24_source_25_idle <= 1;
      end 
      if(_set_flag_508) begin
        _stream_conv2d_24_source_26_source_mode <= 5'b10;
        _stream_conv2d_24_source_26_source_offset <= conv2d_24_stream_act_local_6 + conv2d_24_act_page_comp_offset_buf_2;
      end 
      if(_set_flag_508) begin
        _source_stream_conv2d_24_source_26_pat_size_0 <= cparam_conv2d_24_stream_reduce_size;
        _source_stream_conv2d_24_source_26_pat_stride_0 <= 1;
      end 
      if(_set_flag_508) begin
        _source_stream_conv2d_24_source_26_pat_size_1 <= conv2d_24_next_stream_num_ops;
        _source_stream_conv2d_24_source_26_pat_stride_1 <= 0;
      end 
      if(_set_flag_508) begin
        _source_stream_conv2d_24_source_26_pat_size_2 <= 1;
        _source_stream_conv2d_24_source_26_pat_stride_2 <= 0;
      end 
      if(_set_flag_508) begin
        _source_stream_conv2d_24_source_26_pat_size_3 <= 1;
        _source_stream_conv2d_24_source_26_pat_stride_3 <= 0;
      end 
      if(_set_flag_508) begin
        _stream_conv2d_24_source_26_source_sel <= 9;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_26_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_26_source_offset_buf <= _stream_conv2d_24_source_26_source_offset;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_26_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_26_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_26_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_26_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_26_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_26_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_26_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_26_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_26_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_26_pat_count_0 <= _source_stream_conv2d_24_source_26_pat_size_0 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_26_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_26_pat_count_1 <= _source_stream_conv2d_24_source_26_pat_size_1 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_26_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_26_pat_count_2 <= _source_stream_conv2d_24_source_26_pat_size_2 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_26_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_26_pat_count_3 <= _source_stream_conv2d_24_source_26_pat_size_3 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_26_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_26_pat_size_buf_0 <= _source_stream_conv2d_24_source_26_pat_size_0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_26_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_26_pat_size_buf_1 <= _source_stream_conv2d_24_source_26_pat_size_1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_26_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_26_pat_size_buf_2 <= _source_stream_conv2d_24_source_26_pat_size_2;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_26_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_26_pat_size_buf_3 <= _source_stream_conv2d_24_source_26_pat_size_3;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_26_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_26_pat_stride_buf_0 <= _source_stream_conv2d_24_source_26_pat_stride_0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_26_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_26_pat_stride_buf_1 <= _source_stream_conv2d_24_source_26_pat_stride_1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_26_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_26_pat_stride_buf_2 <= _source_stream_conv2d_24_source_26_pat_stride_2;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_26_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_26_pat_stride_buf_3 <= _source_stream_conv2d_24_source_26_pat_stride_3;
      end 
      if(_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_busy && _stream_conv2d_24_is_root) begin
        __variable_wdata_364 <= _stream_conv2d_24_source_26_source_ram_rdata;
      end 
      if((_stream_conv2d_24_source_26_source_pat_fsm_8 == 1) && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_26_idle <= 0;
        _stream_conv2d_24_source_26_source_ram_raddr <= _stream_conv2d_24_source_26_source_pat_all_offset;
        _stream_conv2d_24_source_26_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_24_source_26_source_pat_fsm_8 == 1) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_26_pat_cur_offset_0 <= _source_stream_conv2d_24_source_26_pat_cur_offset_0 + _source_stream_conv2d_24_source_26_pat_stride_buf_0;
        _source_stream_conv2d_24_source_26_pat_count_0 <= _source_stream_conv2d_24_source_26_pat_count_0 - 1;
      end 
      if((_stream_conv2d_24_source_26_source_pat_fsm_8 == 1) && (_source_stream_conv2d_24_source_26_pat_count_0 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_26_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_24_source_26_pat_count_0 <= _source_stream_conv2d_24_source_26_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_24_source_26_source_pat_fsm_8 == 1) && (_source_stream_conv2d_24_source_26_pat_count_0 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_26_pat_cur_offset_1 <= _source_stream_conv2d_24_source_26_pat_cur_offset_1 + _source_stream_conv2d_24_source_26_pat_stride_buf_1;
        _source_stream_conv2d_24_source_26_pat_count_1 <= _source_stream_conv2d_24_source_26_pat_count_1 - 1;
      end 
      if((_stream_conv2d_24_source_26_source_pat_fsm_8 == 1) && (_source_stream_conv2d_24_source_26_pat_count_0 == 0) && (_source_stream_conv2d_24_source_26_pat_count_1 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_26_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_24_source_26_pat_count_1 <= _source_stream_conv2d_24_source_26_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_24_source_26_source_pat_fsm_8 == 1) && ((_source_stream_conv2d_24_source_26_pat_count_0 == 0) && (_source_stream_conv2d_24_source_26_pat_count_1 == 0)) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_26_pat_cur_offset_2 <= _source_stream_conv2d_24_source_26_pat_cur_offset_2 + _source_stream_conv2d_24_source_26_pat_stride_buf_2;
        _source_stream_conv2d_24_source_26_pat_count_2 <= _source_stream_conv2d_24_source_26_pat_count_2 - 1;
      end 
      if((_stream_conv2d_24_source_26_source_pat_fsm_8 == 1) && ((_source_stream_conv2d_24_source_26_pat_count_0 == 0) && (_source_stream_conv2d_24_source_26_pat_count_1 == 0)) && (_source_stream_conv2d_24_source_26_pat_count_2 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_26_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_24_source_26_pat_count_2 <= _source_stream_conv2d_24_source_26_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_24_source_26_source_pat_fsm_8 == 1) && ((_source_stream_conv2d_24_source_26_pat_count_0 == 0) && (_source_stream_conv2d_24_source_26_pat_count_1 == 0) && (_source_stream_conv2d_24_source_26_pat_count_2 == 0)) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_26_pat_cur_offset_3 <= _source_stream_conv2d_24_source_26_pat_cur_offset_3 + _source_stream_conv2d_24_source_26_pat_stride_buf_3;
        _source_stream_conv2d_24_source_26_pat_count_3 <= _source_stream_conv2d_24_source_26_pat_count_3 - 1;
      end 
      if((_stream_conv2d_24_source_26_source_pat_fsm_8 == 1) && ((_source_stream_conv2d_24_source_26_pat_count_0 == 0) && (_source_stream_conv2d_24_source_26_pat_count_1 == 0) && (_source_stream_conv2d_24_source_26_pat_count_2 == 0)) && (_source_stream_conv2d_24_source_26_pat_count_3 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_26_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_24_source_26_pat_count_3 <= _source_stream_conv2d_24_source_26_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_24_source_26_source_pat_fsm_8 == 1) && _stream_conv2d_24_source_stop && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_26_source_ram_renable <= 0;
        _stream_conv2d_24_source_26_idle <= 1;
      end 
      if((_stream_conv2d_24_source_26_source_pat_fsm_8 == 2) && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_26_source_ram_renable <= 0;
        _stream_conv2d_24_source_26_idle <= 1;
      end 
      if(_set_flag_521) begin
        _stream_conv2d_24_source_27_source_mode <= 5'b10;
        _stream_conv2d_24_source_27_source_offset <= conv2d_24_stream_act_local_7 + conv2d_24_act_page_comp_offset_buf_2;
      end 
      if(_set_flag_521) begin
        _source_stream_conv2d_24_source_27_pat_size_0 <= cparam_conv2d_24_stream_reduce_size;
        _source_stream_conv2d_24_source_27_pat_stride_0 <= 1;
      end 
      if(_set_flag_521) begin
        _source_stream_conv2d_24_source_27_pat_size_1 <= conv2d_24_next_stream_num_ops;
        _source_stream_conv2d_24_source_27_pat_stride_1 <= 0;
      end 
      if(_set_flag_521) begin
        _source_stream_conv2d_24_source_27_pat_size_2 <= 1;
        _source_stream_conv2d_24_source_27_pat_stride_2 <= 0;
      end 
      if(_set_flag_521) begin
        _source_stream_conv2d_24_source_27_pat_size_3 <= 1;
        _source_stream_conv2d_24_source_27_pat_stride_3 <= 0;
      end 
      if(_set_flag_521) begin
        _stream_conv2d_24_source_27_source_sel <= 10;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_27_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_27_source_offset_buf <= _stream_conv2d_24_source_27_source_offset;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_27_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_27_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_27_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_27_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_27_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_27_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_27_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_27_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_27_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_27_pat_count_0 <= _source_stream_conv2d_24_source_27_pat_size_0 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_27_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_27_pat_count_1 <= _source_stream_conv2d_24_source_27_pat_size_1 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_27_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_27_pat_count_2 <= _source_stream_conv2d_24_source_27_pat_size_2 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_27_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_27_pat_count_3 <= _source_stream_conv2d_24_source_27_pat_size_3 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_27_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_27_pat_size_buf_0 <= _source_stream_conv2d_24_source_27_pat_size_0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_27_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_27_pat_size_buf_1 <= _source_stream_conv2d_24_source_27_pat_size_1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_27_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_27_pat_size_buf_2 <= _source_stream_conv2d_24_source_27_pat_size_2;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_27_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_27_pat_size_buf_3 <= _source_stream_conv2d_24_source_27_pat_size_3;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_27_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_27_pat_stride_buf_0 <= _source_stream_conv2d_24_source_27_pat_stride_0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_27_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_27_pat_stride_buf_1 <= _source_stream_conv2d_24_source_27_pat_stride_1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_27_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_27_pat_stride_buf_2 <= _source_stream_conv2d_24_source_27_pat_stride_2;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_27_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_27_pat_stride_buf_3 <= _source_stream_conv2d_24_source_27_pat_stride_3;
      end 
      if(_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_busy && _stream_conv2d_24_is_root) begin
        __variable_wdata_365 <= _stream_conv2d_24_source_27_source_ram_rdata;
      end 
      if((_stream_conv2d_24_source_27_source_pat_fsm_9 == 1) && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_27_idle <= 0;
        _stream_conv2d_24_source_27_source_ram_raddr <= _stream_conv2d_24_source_27_source_pat_all_offset;
        _stream_conv2d_24_source_27_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_24_source_27_source_pat_fsm_9 == 1) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_27_pat_cur_offset_0 <= _source_stream_conv2d_24_source_27_pat_cur_offset_0 + _source_stream_conv2d_24_source_27_pat_stride_buf_0;
        _source_stream_conv2d_24_source_27_pat_count_0 <= _source_stream_conv2d_24_source_27_pat_count_0 - 1;
      end 
      if((_stream_conv2d_24_source_27_source_pat_fsm_9 == 1) && (_source_stream_conv2d_24_source_27_pat_count_0 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_27_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_24_source_27_pat_count_0 <= _source_stream_conv2d_24_source_27_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_24_source_27_source_pat_fsm_9 == 1) && (_source_stream_conv2d_24_source_27_pat_count_0 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_27_pat_cur_offset_1 <= _source_stream_conv2d_24_source_27_pat_cur_offset_1 + _source_stream_conv2d_24_source_27_pat_stride_buf_1;
        _source_stream_conv2d_24_source_27_pat_count_1 <= _source_stream_conv2d_24_source_27_pat_count_1 - 1;
      end 
      if((_stream_conv2d_24_source_27_source_pat_fsm_9 == 1) && (_source_stream_conv2d_24_source_27_pat_count_0 == 0) && (_source_stream_conv2d_24_source_27_pat_count_1 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_27_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_24_source_27_pat_count_1 <= _source_stream_conv2d_24_source_27_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_24_source_27_source_pat_fsm_9 == 1) && ((_source_stream_conv2d_24_source_27_pat_count_0 == 0) && (_source_stream_conv2d_24_source_27_pat_count_1 == 0)) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_27_pat_cur_offset_2 <= _source_stream_conv2d_24_source_27_pat_cur_offset_2 + _source_stream_conv2d_24_source_27_pat_stride_buf_2;
        _source_stream_conv2d_24_source_27_pat_count_2 <= _source_stream_conv2d_24_source_27_pat_count_2 - 1;
      end 
      if((_stream_conv2d_24_source_27_source_pat_fsm_9 == 1) && ((_source_stream_conv2d_24_source_27_pat_count_0 == 0) && (_source_stream_conv2d_24_source_27_pat_count_1 == 0)) && (_source_stream_conv2d_24_source_27_pat_count_2 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_27_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_24_source_27_pat_count_2 <= _source_stream_conv2d_24_source_27_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_24_source_27_source_pat_fsm_9 == 1) && ((_source_stream_conv2d_24_source_27_pat_count_0 == 0) && (_source_stream_conv2d_24_source_27_pat_count_1 == 0) && (_source_stream_conv2d_24_source_27_pat_count_2 == 0)) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_27_pat_cur_offset_3 <= _source_stream_conv2d_24_source_27_pat_cur_offset_3 + _source_stream_conv2d_24_source_27_pat_stride_buf_3;
        _source_stream_conv2d_24_source_27_pat_count_3 <= _source_stream_conv2d_24_source_27_pat_count_3 - 1;
      end 
      if((_stream_conv2d_24_source_27_source_pat_fsm_9 == 1) && ((_source_stream_conv2d_24_source_27_pat_count_0 == 0) && (_source_stream_conv2d_24_source_27_pat_count_1 == 0) && (_source_stream_conv2d_24_source_27_pat_count_2 == 0)) && (_source_stream_conv2d_24_source_27_pat_count_3 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_27_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_24_source_27_pat_count_3 <= _source_stream_conv2d_24_source_27_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_24_source_27_source_pat_fsm_9 == 1) && _stream_conv2d_24_source_stop && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_27_source_ram_renable <= 0;
        _stream_conv2d_24_source_27_idle <= 1;
      end 
      if((_stream_conv2d_24_source_27_source_pat_fsm_9 == 2) && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_27_source_ram_renable <= 0;
        _stream_conv2d_24_source_27_idle <= 1;
      end 
      if(_set_flag_534) begin
        _stream_conv2d_24_source_28_source_mode <= 5'b10;
        _stream_conv2d_24_source_28_source_offset <= conv2d_24_stream_act_local_8 + conv2d_24_act_page_comp_offset_buf_2;
      end 
      if(_set_flag_534) begin
        _source_stream_conv2d_24_source_28_pat_size_0 <= cparam_conv2d_24_stream_reduce_size;
        _source_stream_conv2d_24_source_28_pat_stride_0 <= 1;
      end 
      if(_set_flag_534) begin
        _source_stream_conv2d_24_source_28_pat_size_1 <= conv2d_24_next_stream_num_ops;
        _source_stream_conv2d_24_source_28_pat_stride_1 <= 0;
      end 
      if(_set_flag_534) begin
        _source_stream_conv2d_24_source_28_pat_size_2 <= 1;
        _source_stream_conv2d_24_source_28_pat_stride_2 <= 0;
      end 
      if(_set_flag_534) begin
        _source_stream_conv2d_24_source_28_pat_size_3 <= 1;
        _source_stream_conv2d_24_source_28_pat_stride_3 <= 0;
      end 
      if(_set_flag_534) begin
        _stream_conv2d_24_source_28_source_sel <= 11;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_28_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_28_source_offset_buf <= _stream_conv2d_24_source_28_source_offset;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_28_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_28_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_28_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_28_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_28_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_28_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_28_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_28_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_28_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_28_pat_count_0 <= _source_stream_conv2d_24_source_28_pat_size_0 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_28_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_28_pat_count_1 <= _source_stream_conv2d_24_source_28_pat_size_1 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_28_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_28_pat_count_2 <= _source_stream_conv2d_24_source_28_pat_size_2 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_28_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_28_pat_count_3 <= _source_stream_conv2d_24_source_28_pat_size_3 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_28_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_28_pat_size_buf_0 <= _source_stream_conv2d_24_source_28_pat_size_0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_28_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_28_pat_size_buf_1 <= _source_stream_conv2d_24_source_28_pat_size_1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_28_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_28_pat_size_buf_2 <= _source_stream_conv2d_24_source_28_pat_size_2;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_28_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_28_pat_size_buf_3 <= _source_stream_conv2d_24_source_28_pat_size_3;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_28_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_28_pat_stride_buf_0 <= _source_stream_conv2d_24_source_28_pat_stride_0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_28_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_28_pat_stride_buf_1 <= _source_stream_conv2d_24_source_28_pat_stride_1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_28_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_28_pat_stride_buf_2 <= _source_stream_conv2d_24_source_28_pat_stride_2;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_28_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_28_pat_stride_buf_3 <= _source_stream_conv2d_24_source_28_pat_stride_3;
      end 
      if(_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_busy && _stream_conv2d_24_is_root) begin
        __variable_wdata_366 <= _stream_conv2d_24_source_28_source_ram_rdata;
      end 
      if((_stream_conv2d_24_source_28_source_pat_fsm_10 == 1) && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_28_idle <= 0;
        _stream_conv2d_24_source_28_source_ram_raddr <= _stream_conv2d_24_source_28_source_pat_all_offset;
        _stream_conv2d_24_source_28_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_24_source_28_source_pat_fsm_10 == 1) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_28_pat_cur_offset_0 <= _source_stream_conv2d_24_source_28_pat_cur_offset_0 + _source_stream_conv2d_24_source_28_pat_stride_buf_0;
        _source_stream_conv2d_24_source_28_pat_count_0 <= _source_stream_conv2d_24_source_28_pat_count_0 - 1;
      end 
      if((_stream_conv2d_24_source_28_source_pat_fsm_10 == 1) && (_source_stream_conv2d_24_source_28_pat_count_0 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_28_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_24_source_28_pat_count_0 <= _source_stream_conv2d_24_source_28_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_24_source_28_source_pat_fsm_10 == 1) && (_source_stream_conv2d_24_source_28_pat_count_0 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_28_pat_cur_offset_1 <= _source_stream_conv2d_24_source_28_pat_cur_offset_1 + _source_stream_conv2d_24_source_28_pat_stride_buf_1;
        _source_stream_conv2d_24_source_28_pat_count_1 <= _source_stream_conv2d_24_source_28_pat_count_1 - 1;
      end 
      if((_stream_conv2d_24_source_28_source_pat_fsm_10 == 1) && (_source_stream_conv2d_24_source_28_pat_count_0 == 0) && (_source_stream_conv2d_24_source_28_pat_count_1 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_28_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_24_source_28_pat_count_1 <= _source_stream_conv2d_24_source_28_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_24_source_28_source_pat_fsm_10 == 1) && ((_source_stream_conv2d_24_source_28_pat_count_0 == 0) && (_source_stream_conv2d_24_source_28_pat_count_1 == 0)) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_28_pat_cur_offset_2 <= _source_stream_conv2d_24_source_28_pat_cur_offset_2 + _source_stream_conv2d_24_source_28_pat_stride_buf_2;
        _source_stream_conv2d_24_source_28_pat_count_2 <= _source_stream_conv2d_24_source_28_pat_count_2 - 1;
      end 
      if((_stream_conv2d_24_source_28_source_pat_fsm_10 == 1) && ((_source_stream_conv2d_24_source_28_pat_count_0 == 0) && (_source_stream_conv2d_24_source_28_pat_count_1 == 0)) && (_source_stream_conv2d_24_source_28_pat_count_2 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_28_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_24_source_28_pat_count_2 <= _source_stream_conv2d_24_source_28_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_24_source_28_source_pat_fsm_10 == 1) && ((_source_stream_conv2d_24_source_28_pat_count_0 == 0) && (_source_stream_conv2d_24_source_28_pat_count_1 == 0) && (_source_stream_conv2d_24_source_28_pat_count_2 == 0)) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_28_pat_cur_offset_3 <= _source_stream_conv2d_24_source_28_pat_cur_offset_3 + _source_stream_conv2d_24_source_28_pat_stride_buf_3;
        _source_stream_conv2d_24_source_28_pat_count_3 <= _source_stream_conv2d_24_source_28_pat_count_3 - 1;
      end 
      if((_stream_conv2d_24_source_28_source_pat_fsm_10 == 1) && ((_source_stream_conv2d_24_source_28_pat_count_0 == 0) && (_source_stream_conv2d_24_source_28_pat_count_1 == 0) && (_source_stream_conv2d_24_source_28_pat_count_2 == 0)) && (_source_stream_conv2d_24_source_28_pat_count_3 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_28_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_24_source_28_pat_count_3 <= _source_stream_conv2d_24_source_28_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_24_source_28_source_pat_fsm_10 == 1) && _stream_conv2d_24_source_stop && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_28_source_ram_renable <= 0;
        _stream_conv2d_24_source_28_idle <= 1;
      end 
      if((_stream_conv2d_24_source_28_source_pat_fsm_10 == 2) && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_28_source_ram_renable <= 0;
        _stream_conv2d_24_source_28_idle <= 1;
      end 
      if(_set_flag_547) begin
        _stream_conv2d_24_source_29_source_mode <= 5'b10;
        _stream_conv2d_24_source_29_source_offset <= conv2d_24_filter_page_comp_offset_buf;
      end 
      if(_set_flag_547) begin
        _source_stream_conv2d_24_source_29_pat_size_0 <= cparam_conv2d_24_stream_reduce_size;
        _source_stream_conv2d_24_source_29_pat_stride_0 <= 1;
      end 
      if(_set_flag_547) begin
        _source_stream_conv2d_24_source_29_pat_size_1 <= conv2d_24_next_stream_num_ops;
        _source_stream_conv2d_24_source_29_pat_stride_1 <= cparam_conv2d_24_stream_aligned_reduce_size;
      end 
      if(_set_flag_547) begin
        _source_stream_conv2d_24_source_29_pat_size_2 <= 1;
        _source_stream_conv2d_24_source_29_pat_stride_2 <= 0;
      end 
      if(_set_flag_547) begin
        _source_stream_conv2d_24_source_29_pat_size_3 <= 1;
        _source_stream_conv2d_24_source_29_pat_stride_3 <= 0;
      end 
      if(_set_flag_547) begin
        _stream_conv2d_24_source_29_source_sel <= 12;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_29_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_29_source_offset_buf <= _stream_conv2d_24_source_29_source_offset;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_29_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_29_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_29_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_29_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_29_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_29_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_29_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_29_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_29_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_29_pat_count_0 <= _source_stream_conv2d_24_source_29_pat_size_0 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_29_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_29_pat_count_1 <= _source_stream_conv2d_24_source_29_pat_size_1 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_29_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_29_pat_count_2 <= _source_stream_conv2d_24_source_29_pat_size_2 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_29_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_29_pat_count_3 <= _source_stream_conv2d_24_source_29_pat_size_3 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_29_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_29_pat_size_buf_0 <= _source_stream_conv2d_24_source_29_pat_size_0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_29_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_29_pat_size_buf_1 <= _source_stream_conv2d_24_source_29_pat_size_1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_29_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_29_pat_size_buf_2 <= _source_stream_conv2d_24_source_29_pat_size_2;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_29_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_29_pat_size_buf_3 <= _source_stream_conv2d_24_source_29_pat_size_3;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_29_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_29_pat_stride_buf_0 <= _source_stream_conv2d_24_source_29_pat_stride_0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_29_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_29_pat_stride_buf_1 <= _source_stream_conv2d_24_source_29_pat_stride_1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_29_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_29_pat_stride_buf_2 <= _source_stream_conv2d_24_source_29_pat_stride_2;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_29_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_29_pat_stride_buf_3 <= _source_stream_conv2d_24_source_29_pat_stride_3;
      end 
      if(_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_busy && _stream_conv2d_24_is_root) begin
        __variable_wdata_592 <= _stream_conv2d_24_source_29_source_ram_rdata;
      end 
      if((_stream_conv2d_24_source_29_source_pat_fsm_11 == 1) && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_29_idle <= 0;
        _stream_conv2d_24_source_29_source_ram_raddr <= _stream_conv2d_24_source_29_source_pat_all_offset;
        _stream_conv2d_24_source_29_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_24_source_29_source_pat_fsm_11 == 1) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_29_pat_cur_offset_0 <= _source_stream_conv2d_24_source_29_pat_cur_offset_0 + _source_stream_conv2d_24_source_29_pat_stride_buf_0;
        _source_stream_conv2d_24_source_29_pat_count_0 <= _source_stream_conv2d_24_source_29_pat_count_0 - 1;
      end 
      if((_stream_conv2d_24_source_29_source_pat_fsm_11 == 1) && (_source_stream_conv2d_24_source_29_pat_count_0 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_29_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_24_source_29_pat_count_0 <= _source_stream_conv2d_24_source_29_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_24_source_29_source_pat_fsm_11 == 1) && (_source_stream_conv2d_24_source_29_pat_count_0 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_29_pat_cur_offset_1 <= _source_stream_conv2d_24_source_29_pat_cur_offset_1 + _source_stream_conv2d_24_source_29_pat_stride_buf_1;
        _source_stream_conv2d_24_source_29_pat_count_1 <= _source_stream_conv2d_24_source_29_pat_count_1 - 1;
      end 
      if((_stream_conv2d_24_source_29_source_pat_fsm_11 == 1) && (_source_stream_conv2d_24_source_29_pat_count_0 == 0) && (_source_stream_conv2d_24_source_29_pat_count_1 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_29_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_24_source_29_pat_count_1 <= _source_stream_conv2d_24_source_29_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_24_source_29_source_pat_fsm_11 == 1) && ((_source_stream_conv2d_24_source_29_pat_count_0 == 0) && (_source_stream_conv2d_24_source_29_pat_count_1 == 0)) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_29_pat_cur_offset_2 <= _source_stream_conv2d_24_source_29_pat_cur_offset_2 + _source_stream_conv2d_24_source_29_pat_stride_buf_2;
        _source_stream_conv2d_24_source_29_pat_count_2 <= _source_stream_conv2d_24_source_29_pat_count_2 - 1;
      end 
      if((_stream_conv2d_24_source_29_source_pat_fsm_11 == 1) && ((_source_stream_conv2d_24_source_29_pat_count_0 == 0) && (_source_stream_conv2d_24_source_29_pat_count_1 == 0)) && (_source_stream_conv2d_24_source_29_pat_count_2 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_29_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_24_source_29_pat_count_2 <= _source_stream_conv2d_24_source_29_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_24_source_29_source_pat_fsm_11 == 1) && ((_source_stream_conv2d_24_source_29_pat_count_0 == 0) && (_source_stream_conv2d_24_source_29_pat_count_1 == 0) && (_source_stream_conv2d_24_source_29_pat_count_2 == 0)) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_29_pat_cur_offset_3 <= _source_stream_conv2d_24_source_29_pat_cur_offset_3 + _source_stream_conv2d_24_source_29_pat_stride_buf_3;
        _source_stream_conv2d_24_source_29_pat_count_3 <= _source_stream_conv2d_24_source_29_pat_count_3 - 1;
      end 
      if((_stream_conv2d_24_source_29_source_pat_fsm_11 == 1) && ((_source_stream_conv2d_24_source_29_pat_count_0 == 0) && (_source_stream_conv2d_24_source_29_pat_count_1 == 0) && (_source_stream_conv2d_24_source_29_pat_count_2 == 0)) && (_source_stream_conv2d_24_source_29_pat_count_3 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_29_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_24_source_29_pat_count_3 <= _source_stream_conv2d_24_source_29_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_24_source_29_source_pat_fsm_11 == 1) && _stream_conv2d_24_source_stop && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_29_source_ram_renable <= 0;
        _stream_conv2d_24_source_29_idle <= 1;
      end 
      if((_stream_conv2d_24_source_29_source_pat_fsm_11 == 2) && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_29_source_ram_renable <= 0;
        _stream_conv2d_24_source_29_idle <= 1;
      end 
      if(_set_flag_560) begin
        _stream_conv2d_24_source_30_source_mode <= 5'b10;
        _stream_conv2d_24_source_30_source_offset <= conv2d_24_filter_page_comp_offset_buf;
      end 
      if(_set_flag_560) begin
        _source_stream_conv2d_24_source_30_pat_size_0 <= cparam_conv2d_24_stream_reduce_size;
        _source_stream_conv2d_24_source_30_pat_stride_0 <= 1;
      end 
      if(_set_flag_560) begin
        _source_stream_conv2d_24_source_30_pat_size_1 <= conv2d_24_next_stream_num_ops;
        _source_stream_conv2d_24_source_30_pat_stride_1 <= cparam_conv2d_24_stream_aligned_reduce_size;
      end 
      if(_set_flag_560) begin
        _source_stream_conv2d_24_source_30_pat_size_2 <= 1;
        _source_stream_conv2d_24_source_30_pat_stride_2 <= 0;
      end 
      if(_set_flag_560) begin
        _source_stream_conv2d_24_source_30_pat_size_3 <= 1;
        _source_stream_conv2d_24_source_30_pat_stride_3 <= 0;
      end 
      if(_set_flag_560) begin
        _stream_conv2d_24_source_30_source_sel <= 13;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_30_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_30_source_offset_buf <= _stream_conv2d_24_source_30_source_offset;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_30_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_30_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_30_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_30_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_30_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_30_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_30_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_30_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_30_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_30_pat_count_0 <= _source_stream_conv2d_24_source_30_pat_size_0 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_30_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_30_pat_count_1 <= _source_stream_conv2d_24_source_30_pat_size_1 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_30_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_30_pat_count_2 <= _source_stream_conv2d_24_source_30_pat_size_2 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_30_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_30_pat_count_3 <= _source_stream_conv2d_24_source_30_pat_size_3 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_30_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_30_pat_size_buf_0 <= _source_stream_conv2d_24_source_30_pat_size_0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_30_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_30_pat_size_buf_1 <= _source_stream_conv2d_24_source_30_pat_size_1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_30_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_30_pat_size_buf_2 <= _source_stream_conv2d_24_source_30_pat_size_2;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_30_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_30_pat_size_buf_3 <= _source_stream_conv2d_24_source_30_pat_size_3;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_30_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_30_pat_stride_buf_0 <= _source_stream_conv2d_24_source_30_pat_stride_0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_30_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_30_pat_stride_buf_1 <= _source_stream_conv2d_24_source_30_pat_stride_1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_30_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_30_pat_stride_buf_2 <= _source_stream_conv2d_24_source_30_pat_stride_2;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_30_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_30_pat_stride_buf_3 <= _source_stream_conv2d_24_source_30_pat_stride_3;
      end 
      if(_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_busy && _stream_conv2d_24_is_root) begin
        __variable_wdata_593 <= _stream_conv2d_24_source_30_source_ram_rdata;
      end 
      if((_stream_conv2d_24_source_30_source_pat_fsm_12 == 1) && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_30_idle <= 0;
        _stream_conv2d_24_source_30_source_ram_raddr <= _stream_conv2d_24_source_30_source_pat_all_offset;
        _stream_conv2d_24_source_30_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_24_source_30_source_pat_fsm_12 == 1) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_30_pat_cur_offset_0 <= _source_stream_conv2d_24_source_30_pat_cur_offset_0 + _source_stream_conv2d_24_source_30_pat_stride_buf_0;
        _source_stream_conv2d_24_source_30_pat_count_0 <= _source_stream_conv2d_24_source_30_pat_count_0 - 1;
      end 
      if((_stream_conv2d_24_source_30_source_pat_fsm_12 == 1) && (_source_stream_conv2d_24_source_30_pat_count_0 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_30_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_24_source_30_pat_count_0 <= _source_stream_conv2d_24_source_30_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_24_source_30_source_pat_fsm_12 == 1) && (_source_stream_conv2d_24_source_30_pat_count_0 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_30_pat_cur_offset_1 <= _source_stream_conv2d_24_source_30_pat_cur_offset_1 + _source_stream_conv2d_24_source_30_pat_stride_buf_1;
        _source_stream_conv2d_24_source_30_pat_count_1 <= _source_stream_conv2d_24_source_30_pat_count_1 - 1;
      end 
      if((_stream_conv2d_24_source_30_source_pat_fsm_12 == 1) && (_source_stream_conv2d_24_source_30_pat_count_0 == 0) && (_source_stream_conv2d_24_source_30_pat_count_1 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_30_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_24_source_30_pat_count_1 <= _source_stream_conv2d_24_source_30_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_24_source_30_source_pat_fsm_12 == 1) && ((_source_stream_conv2d_24_source_30_pat_count_0 == 0) && (_source_stream_conv2d_24_source_30_pat_count_1 == 0)) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_30_pat_cur_offset_2 <= _source_stream_conv2d_24_source_30_pat_cur_offset_2 + _source_stream_conv2d_24_source_30_pat_stride_buf_2;
        _source_stream_conv2d_24_source_30_pat_count_2 <= _source_stream_conv2d_24_source_30_pat_count_2 - 1;
      end 
      if((_stream_conv2d_24_source_30_source_pat_fsm_12 == 1) && ((_source_stream_conv2d_24_source_30_pat_count_0 == 0) && (_source_stream_conv2d_24_source_30_pat_count_1 == 0)) && (_source_stream_conv2d_24_source_30_pat_count_2 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_30_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_24_source_30_pat_count_2 <= _source_stream_conv2d_24_source_30_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_24_source_30_source_pat_fsm_12 == 1) && ((_source_stream_conv2d_24_source_30_pat_count_0 == 0) && (_source_stream_conv2d_24_source_30_pat_count_1 == 0) && (_source_stream_conv2d_24_source_30_pat_count_2 == 0)) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_30_pat_cur_offset_3 <= _source_stream_conv2d_24_source_30_pat_cur_offset_3 + _source_stream_conv2d_24_source_30_pat_stride_buf_3;
        _source_stream_conv2d_24_source_30_pat_count_3 <= _source_stream_conv2d_24_source_30_pat_count_3 - 1;
      end 
      if((_stream_conv2d_24_source_30_source_pat_fsm_12 == 1) && ((_source_stream_conv2d_24_source_30_pat_count_0 == 0) && (_source_stream_conv2d_24_source_30_pat_count_1 == 0) && (_source_stream_conv2d_24_source_30_pat_count_2 == 0)) && (_source_stream_conv2d_24_source_30_pat_count_3 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_30_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_24_source_30_pat_count_3 <= _source_stream_conv2d_24_source_30_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_24_source_30_source_pat_fsm_12 == 1) && _stream_conv2d_24_source_stop && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_30_source_ram_renable <= 0;
        _stream_conv2d_24_source_30_idle <= 1;
      end 
      if((_stream_conv2d_24_source_30_source_pat_fsm_12 == 2) && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_30_source_ram_renable <= 0;
        _stream_conv2d_24_source_30_idle <= 1;
      end 
      if(_set_flag_573) begin
        _stream_conv2d_24_source_31_source_mode <= 5'b10;
        _stream_conv2d_24_source_31_source_offset <= conv2d_24_filter_page_comp_offset_buf;
      end 
      if(_set_flag_573) begin
        _source_stream_conv2d_24_source_31_pat_size_0 <= cparam_conv2d_24_stream_reduce_size;
        _source_stream_conv2d_24_source_31_pat_stride_0 <= 1;
      end 
      if(_set_flag_573) begin
        _source_stream_conv2d_24_source_31_pat_size_1 <= conv2d_24_next_stream_num_ops;
        _source_stream_conv2d_24_source_31_pat_stride_1 <= cparam_conv2d_24_stream_aligned_reduce_size;
      end 
      if(_set_flag_573) begin
        _source_stream_conv2d_24_source_31_pat_size_2 <= 1;
        _source_stream_conv2d_24_source_31_pat_stride_2 <= 0;
      end 
      if(_set_flag_573) begin
        _source_stream_conv2d_24_source_31_pat_size_3 <= 1;
        _source_stream_conv2d_24_source_31_pat_stride_3 <= 0;
      end 
      if(_set_flag_573) begin
        _stream_conv2d_24_source_31_source_sel <= 14;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_31_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_31_source_offset_buf <= _stream_conv2d_24_source_31_source_offset;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_31_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_31_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_31_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_31_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_31_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_31_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_31_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_31_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_31_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_31_pat_count_0 <= _source_stream_conv2d_24_source_31_pat_size_0 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_31_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_31_pat_count_1 <= _source_stream_conv2d_24_source_31_pat_size_1 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_31_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_31_pat_count_2 <= _source_stream_conv2d_24_source_31_pat_size_2 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_31_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_31_pat_count_3 <= _source_stream_conv2d_24_source_31_pat_size_3 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_31_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_31_pat_size_buf_0 <= _source_stream_conv2d_24_source_31_pat_size_0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_31_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_31_pat_size_buf_1 <= _source_stream_conv2d_24_source_31_pat_size_1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_31_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_31_pat_size_buf_2 <= _source_stream_conv2d_24_source_31_pat_size_2;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_31_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_31_pat_size_buf_3 <= _source_stream_conv2d_24_source_31_pat_size_3;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_31_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_31_pat_stride_buf_0 <= _source_stream_conv2d_24_source_31_pat_stride_0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_31_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_31_pat_stride_buf_1 <= _source_stream_conv2d_24_source_31_pat_stride_1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_31_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_31_pat_stride_buf_2 <= _source_stream_conv2d_24_source_31_pat_stride_2;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_31_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_31_pat_stride_buf_3 <= _source_stream_conv2d_24_source_31_pat_stride_3;
      end 
      if(_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_busy && _stream_conv2d_24_is_root) begin
        __variable_wdata_594 <= _stream_conv2d_24_source_31_source_ram_rdata;
      end 
      if((_stream_conv2d_24_source_31_source_pat_fsm_13 == 1) && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_31_idle <= 0;
        _stream_conv2d_24_source_31_source_ram_raddr <= _stream_conv2d_24_source_31_source_pat_all_offset;
        _stream_conv2d_24_source_31_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_24_source_31_source_pat_fsm_13 == 1) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_31_pat_cur_offset_0 <= _source_stream_conv2d_24_source_31_pat_cur_offset_0 + _source_stream_conv2d_24_source_31_pat_stride_buf_0;
        _source_stream_conv2d_24_source_31_pat_count_0 <= _source_stream_conv2d_24_source_31_pat_count_0 - 1;
      end 
      if((_stream_conv2d_24_source_31_source_pat_fsm_13 == 1) && (_source_stream_conv2d_24_source_31_pat_count_0 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_31_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_24_source_31_pat_count_0 <= _source_stream_conv2d_24_source_31_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_24_source_31_source_pat_fsm_13 == 1) && (_source_stream_conv2d_24_source_31_pat_count_0 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_31_pat_cur_offset_1 <= _source_stream_conv2d_24_source_31_pat_cur_offset_1 + _source_stream_conv2d_24_source_31_pat_stride_buf_1;
        _source_stream_conv2d_24_source_31_pat_count_1 <= _source_stream_conv2d_24_source_31_pat_count_1 - 1;
      end 
      if((_stream_conv2d_24_source_31_source_pat_fsm_13 == 1) && (_source_stream_conv2d_24_source_31_pat_count_0 == 0) && (_source_stream_conv2d_24_source_31_pat_count_1 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_31_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_24_source_31_pat_count_1 <= _source_stream_conv2d_24_source_31_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_24_source_31_source_pat_fsm_13 == 1) && ((_source_stream_conv2d_24_source_31_pat_count_0 == 0) && (_source_stream_conv2d_24_source_31_pat_count_1 == 0)) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_31_pat_cur_offset_2 <= _source_stream_conv2d_24_source_31_pat_cur_offset_2 + _source_stream_conv2d_24_source_31_pat_stride_buf_2;
        _source_stream_conv2d_24_source_31_pat_count_2 <= _source_stream_conv2d_24_source_31_pat_count_2 - 1;
      end 
      if((_stream_conv2d_24_source_31_source_pat_fsm_13 == 1) && ((_source_stream_conv2d_24_source_31_pat_count_0 == 0) && (_source_stream_conv2d_24_source_31_pat_count_1 == 0)) && (_source_stream_conv2d_24_source_31_pat_count_2 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_31_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_24_source_31_pat_count_2 <= _source_stream_conv2d_24_source_31_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_24_source_31_source_pat_fsm_13 == 1) && ((_source_stream_conv2d_24_source_31_pat_count_0 == 0) && (_source_stream_conv2d_24_source_31_pat_count_1 == 0) && (_source_stream_conv2d_24_source_31_pat_count_2 == 0)) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_31_pat_cur_offset_3 <= _source_stream_conv2d_24_source_31_pat_cur_offset_3 + _source_stream_conv2d_24_source_31_pat_stride_buf_3;
        _source_stream_conv2d_24_source_31_pat_count_3 <= _source_stream_conv2d_24_source_31_pat_count_3 - 1;
      end 
      if((_stream_conv2d_24_source_31_source_pat_fsm_13 == 1) && ((_source_stream_conv2d_24_source_31_pat_count_0 == 0) && (_source_stream_conv2d_24_source_31_pat_count_1 == 0) && (_source_stream_conv2d_24_source_31_pat_count_2 == 0)) && (_source_stream_conv2d_24_source_31_pat_count_3 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_31_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_24_source_31_pat_count_3 <= _source_stream_conv2d_24_source_31_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_24_source_31_source_pat_fsm_13 == 1) && _stream_conv2d_24_source_stop && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_31_source_ram_renable <= 0;
        _stream_conv2d_24_source_31_idle <= 1;
      end 
      if((_stream_conv2d_24_source_31_source_pat_fsm_13 == 2) && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_31_source_ram_renable <= 0;
        _stream_conv2d_24_source_31_idle <= 1;
      end 
      if(_set_flag_586) begin
        _stream_conv2d_24_source_32_source_mode <= 5'b10;
        _stream_conv2d_24_source_32_source_offset <= conv2d_24_filter_page_comp_offset_buf;
      end 
      if(_set_flag_586) begin
        _source_stream_conv2d_24_source_32_pat_size_0 <= cparam_conv2d_24_stream_reduce_size;
        _source_stream_conv2d_24_source_32_pat_stride_0 <= 1;
      end 
      if(_set_flag_586) begin
        _source_stream_conv2d_24_source_32_pat_size_1 <= conv2d_24_next_stream_num_ops;
        _source_stream_conv2d_24_source_32_pat_stride_1 <= cparam_conv2d_24_stream_aligned_reduce_size;
      end 
      if(_set_flag_586) begin
        _source_stream_conv2d_24_source_32_pat_size_2 <= 1;
        _source_stream_conv2d_24_source_32_pat_stride_2 <= 0;
      end 
      if(_set_flag_586) begin
        _source_stream_conv2d_24_source_32_pat_size_3 <= 1;
        _source_stream_conv2d_24_source_32_pat_stride_3 <= 0;
      end 
      if(_set_flag_586) begin
        _stream_conv2d_24_source_32_source_sel <= 15;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_32_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_32_source_offset_buf <= _stream_conv2d_24_source_32_source_offset;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_32_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_32_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_32_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_32_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_32_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_32_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_32_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_32_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_32_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_32_pat_count_0 <= _source_stream_conv2d_24_source_32_pat_size_0 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_32_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_32_pat_count_1 <= _source_stream_conv2d_24_source_32_pat_size_1 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_32_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_32_pat_count_2 <= _source_stream_conv2d_24_source_32_pat_size_2 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_32_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_32_pat_count_3 <= _source_stream_conv2d_24_source_32_pat_size_3 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_32_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_32_pat_size_buf_0 <= _source_stream_conv2d_24_source_32_pat_size_0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_32_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_32_pat_size_buf_1 <= _source_stream_conv2d_24_source_32_pat_size_1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_32_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_32_pat_size_buf_2 <= _source_stream_conv2d_24_source_32_pat_size_2;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_32_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_32_pat_size_buf_3 <= _source_stream_conv2d_24_source_32_pat_size_3;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_32_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_32_pat_stride_buf_0 <= _source_stream_conv2d_24_source_32_pat_stride_0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_32_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_32_pat_stride_buf_1 <= _source_stream_conv2d_24_source_32_pat_stride_1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_32_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_32_pat_stride_buf_2 <= _source_stream_conv2d_24_source_32_pat_stride_2;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_32_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_32_pat_stride_buf_3 <= _source_stream_conv2d_24_source_32_pat_stride_3;
      end 
      if(_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_busy && _stream_conv2d_24_is_root) begin
        __variable_wdata_595 <= _stream_conv2d_24_source_32_source_ram_rdata;
      end 
      if((_stream_conv2d_24_source_32_source_pat_fsm_14 == 1) && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_32_idle <= 0;
        _stream_conv2d_24_source_32_source_ram_raddr <= _stream_conv2d_24_source_32_source_pat_all_offset;
        _stream_conv2d_24_source_32_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_24_source_32_source_pat_fsm_14 == 1) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_32_pat_cur_offset_0 <= _source_stream_conv2d_24_source_32_pat_cur_offset_0 + _source_stream_conv2d_24_source_32_pat_stride_buf_0;
        _source_stream_conv2d_24_source_32_pat_count_0 <= _source_stream_conv2d_24_source_32_pat_count_0 - 1;
      end 
      if((_stream_conv2d_24_source_32_source_pat_fsm_14 == 1) && (_source_stream_conv2d_24_source_32_pat_count_0 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_32_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_24_source_32_pat_count_0 <= _source_stream_conv2d_24_source_32_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_24_source_32_source_pat_fsm_14 == 1) && (_source_stream_conv2d_24_source_32_pat_count_0 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_32_pat_cur_offset_1 <= _source_stream_conv2d_24_source_32_pat_cur_offset_1 + _source_stream_conv2d_24_source_32_pat_stride_buf_1;
        _source_stream_conv2d_24_source_32_pat_count_1 <= _source_stream_conv2d_24_source_32_pat_count_1 - 1;
      end 
      if((_stream_conv2d_24_source_32_source_pat_fsm_14 == 1) && (_source_stream_conv2d_24_source_32_pat_count_0 == 0) && (_source_stream_conv2d_24_source_32_pat_count_1 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_32_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_24_source_32_pat_count_1 <= _source_stream_conv2d_24_source_32_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_24_source_32_source_pat_fsm_14 == 1) && ((_source_stream_conv2d_24_source_32_pat_count_0 == 0) && (_source_stream_conv2d_24_source_32_pat_count_1 == 0)) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_32_pat_cur_offset_2 <= _source_stream_conv2d_24_source_32_pat_cur_offset_2 + _source_stream_conv2d_24_source_32_pat_stride_buf_2;
        _source_stream_conv2d_24_source_32_pat_count_2 <= _source_stream_conv2d_24_source_32_pat_count_2 - 1;
      end 
      if((_stream_conv2d_24_source_32_source_pat_fsm_14 == 1) && ((_source_stream_conv2d_24_source_32_pat_count_0 == 0) && (_source_stream_conv2d_24_source_32_pat_count_1 == 0)) && (_source_stream_conv2d_24_source_32_pat_count_2 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_32_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_24_source_32_pat_count_2 <= _source_stream_conv2d_24_source_32_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_24_source_32_source_pat_fsm_14 == 1) && ((_source_stream_conv2d_24_source_32_pat_count_0 == 0) && (_source_stream_conv2d_24_source_32_pat_count_1 == 0) && (_source_stream_conv2d_24_source_32_pat_count_2 == 0)) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_32_pat_cur_offset_3 <= _source_stream_conv2d_24_source_32_pat_cur_offset_3 + _source_stream_conv2d_24_source_32_pat_stride_buf_3;
        _source_stream_conv2d_24_source_32_pat_count_3 <= _source_stream_conv2d_24_source_32_pat_count_3 - 1;
      end 
      if((_stream_conv2d_24_source_32_source_pat_fsm_14 == 1) && ((_source_stream_conv2d_24_source_32_pat_count_0 == 0) && (_source_stream_conv2d_24_source_32_pat_count_1 == 0) && (_source_stream_conv2d_24_source_32_pat_count_2 == 0)) && (_source_stream_conv2d_24_source_32_pat_count_3 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_32_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_24_source_32_pat_count_3 <= _source_stream_conv2d_24_source_32_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_24_source_32_source_pat_fsm_14 == 1) && _stream_conv2d_24_source_stop && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_32_source_ram_renable <= 0;
        _stream_conv2d_24_source_32_idle <= 1;
      end 
      if((_stream_conv2d_24_source_32_source_pat_fsm_14 == 2) && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_32_source_ram_renable <= 0;
        _stream_conv2d_24_source_32_idle <= 1;
      end 
      if(_set_flag_599) begin
        _stream_conv2d_24_source_33_source_mode <= 5'b10;
        _stream_conv2d_24_source_33_source_offset <= conv2d_24_filter_page_comp_offset_buf;
      end 
      if(_set_flag_599) begin
        _source_stream_conv2d_24_source_33_pat_size_0 <= cparam_conv2d_24_stream_reduce_size;
        _source_stream_conv2d_24_source_33_pat_stride_0 <= 1;
      end 
      if(_set_flag_599) begin
        _source_stream_conv2d_24_source_33_pat_size_1 <= conv2d_24_next_stream_num_ops;
        _source_stream_conv2d_24_source_33_pat_stride_1 <= cparam_conv2d_24_stream_aligned_reduce_size;
      end 
      if(_set_flag_599) begin
        _source_stream_conv2d_24_source_33_pat_size_2 <= 1;
        _source_stream_conv2d_24_source_33_pat_stride_2 <= 0;
      end 
      if(_set_flag_599) begin
        _source_stream_conv2d_24_source_33_pat_size_3 <= 1;
        _source_stream_conv2d_24_source_33_pat_stride_3 <= 0;
      end 
      if(_set_flag_599) begin
        _stream_conv2d_24_source_33_source_sel <= 16;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_33_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_33_source_offset_buf <= _stream_conv2d_24_source_33_source_offset;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_33_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_33_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_33_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_33_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_33_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_33_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_33_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_33_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_33_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_33_pat_count_0 <= _source_stream_conv2d_24_source_33_pat_size_0 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_33_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_33_pat_count_1 <= _source_stream_conv2d_24_source_33_pat_size_1 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_33_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_33_pat_count_2 <= _source_stream_conv2d_24_source_33_pat_size_2 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_33_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_33_pat_count_3 <= _source_stream_conv2d_24_source_33_pat_size_3 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_33_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_33_pat_size_buf_0 <= _source_stream_conv2d_24_source_33_pat_size_0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_33_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_33_pat_size_buf_1 <= _source_stream_conv2d_24_source_33_pat_size_1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_33_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_33_pat_size_buf_2 <= _source_stream_conv2d_24_source_33_pat_size_2;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_33_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_33_pat_size_buf_3 <= _source_stream_conv2d_24_source_33_pat_size_3;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_33_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_33_pat_stride_buf_0 <= _source_stream_conv2d_24_source_33_pat_stride_0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_33_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_33_pat_stride_buf_1 <= _source_stream_conv2d_24_source_33_pat_stride_1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_33_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_33_pat_stride_buf_2 <= _source_stream_conv2d_24_source_33_pat_stride_2;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_33_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_33_pat_stride_buf_3 <= _source_stream_conv2d_24_source_33_pat_stride_3;
      end 
      if(_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_busy && _stream_conv2d_24_is_root) begin
        __variable_wdata_596 <= _stream_conv2d_24_source_33_source_ram_rdata;
      end 
      if((_stream_conv2d_24_source_33_source_pat_fsm_15 == 1) && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_33_idle <= 0;
        _stream_conv2d_24_source_33_source_ram_raddr <= _stream_conv2d_24_source_33_source_pat_all_offset;
        _stream_conv2d_24_source_33_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_24_source_33_source_pat_fsm_15 == 1) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_33_pat_cur_offset_0 <= _source_stream_conv2d_24_source_33_pat_cur_offset_0 + _source_stream_conv2d_24_source_33_pat_stride_buf_0;
        _source_stream_conv2d_24_source_33_pat_count_0 <= _source_stream_conv2d_24_source_33_pat_count_0 - 1;
      end 
      if((_stream_conv2d_24_source_33_source_pat_fsm_15 == 1) && (_source_stream_conv2d_24_source_33_pat_count_0 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_33_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_24_source_33_pat_count_0 <= _source_stream_conv2d_24_source_33_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_24_source_33_source_pat_fsm_15 == 1) && (_source_stream_conv2d_24_source_33_pat_count_0 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_33_pat_cur_offset_1 <= _source_stream_conv2d_24_source_33_pat_cur_offset_1 + _source_stream_conv2d_24_source_33_pat_stride_buf_1;
        _source_stream_conv2d_24_source_33_pat_count_1 <= _source_stream_conv2d_24_source_33_pat_count_1 - 1;
      end 
      if((_stream_conv2d_24_source_33_source_pat_fsm_15 == 1) && (_source_stream_conv2d_24_source_33_pat_count_0 == 0) && (_source_stream_conv2d_24_source_33_pat_count_1 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_33_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_24_source_33_pat_count_1 <= _source_stream_conv2d_24_source_33_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_24_source_33_source_pat_fsm_15 == 1) && ((_source_stream_conv2d_24_source_33_pat_count_0 == 0) && (_source_stream_conv2d_24_source_33_pat_count_1 == 0)) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_33_pat_cur_offset_2 <= _source_stream_conv2d_24_source_33_pat_cur_offset_2 + _source_stream_conv2d_24_source_33_pat_stride_buf_2;
        _source_stream_conv2d_24_source_33_pat_count_2 <= _source_stream_conv2d_24_source_33_pat_count_2 - 1;
      end 
      if((_stream_conv2d_24_source_33_source_pat_fsm_15 == 1) && ((_source_stream_conv2d_24_source_33_pat_count_0 == 0) && (_source_stream_conv2d_24_source_33_pat_count_1 == 0)) && (_source_stream_conv2d_24_source_33_pat_count_2 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_33_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_24_source_33_pat_count_2 <= _source_stream_conv2d_24_source_33_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_24_source_33_source_pat_fsm_15 == 1) && ((_source_stream_conv2d_24_source_33_pat_count_0 == 0) && (_source_stream_conv2d_24_source_33_pat_count_1 == 0) && (_source_stream_conv2d_24_source_33_pat_count_2 == 0)) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_33_pat_cur_offset_3 <= _source_stream_conv2d_24_source_33_pat_cur_offset_3 + _source_stream_conv2d_24_source_33_pat_stride_buf_3;
        _source_stream_conv2d_24_source_33_pat_count_3 <= _source_stream_conv2d_24_source_33_pat_count_3 - 1;
      end 
      if((_stream_conv2d_24_source_33_source_pat_fsm_15 == 1) && ((_source_stream_conv2d_24_source_33_pat_count_0 == 0) && (_source_stream_conv2d_24_source_33_pat_count_1 == 0) && (_source_stream_conv2d_24_source_33_pat_count_2 == 0)) && (_source_stream_conv2d_24_source_33_pat_count_3 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_33_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_24_source_33_pat_count_3 <= _source_stream_conv2d_24_source_33_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_24_source_33_source_pat_fsm_15 == 1) && _stream_conv2d_24_source_stop && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_33_source_ram_renable <= 0;
        _stream_conv2d_24_source_33_idle <= 1;
      end 
      if((_stream_conv2d_24_source_33_source_pat_fsm_15 == 2) && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_33_source_ram_renable <= 0;
        _stream_conv2d_24_source_33_idle <= 1;
      end 
      if(_set_flag_612) begin
        _stream_conv2d_24_source_34_source_mode <= 5'b10;
        _stream_conv2d_24_source_34_source_offset <= conv2d_24_filter_page_comp_offset_buf;
      end 
      if(_set_flag_612) begin
        _source_stream_conv2d_24_source_34_pat_size_0 <= cparam_conv2d_24_stream_reduce_size;
        _source_stream_conv2d_24_source_34_pat_stride_0 <= 1;
      end 
      if(_set_flag_612) begin
        _source_stream_conv2d_24_source_34_pat_size_1 <= conv2d_24_next_stream_num_ops;
        _source_stream_conv2d_24_source_34_pat_stride_1 <= cparam_conv2d_24_stream_aligned_reduce_size;
      end 
      if(_set_flag_612) begin
        _source_stream_conv2d_24_source_34_pat_size_2 <= 1;
        _source_stream_conv2d_24_source_34_pat_stride_2 <= 0;
      end 
      if(_set_flag_612) begin
        _source_stream_conv2d_24_source_34_pat_size_3 <= 1;
        _source_stream_conv2d_24_source_34_pat_stride_3 <= 0;
      end 
      if(_set_flag_612) begin
        _stream_conv2d_24_source_34_source_sel <= 17;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_34_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_34_source_offset_buf <= _stream_conv2d_24_source_34_source_offset;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_34_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_34_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_34_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_34_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_34_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_34_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_34_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_34_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_34_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_34_pat_count_0 <= _source_stream_conv2d_24_source_34_pat_size_0 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_34_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_34_pat_count_1 <= _source_stream_conv2d_24_source_34_pat_size_1 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_34_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_34_pat_count_2 <= _source_stream_conv2d_24_source_34_pat_size_2 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_34_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_34_pat_count_3 <= _source_stream_conv2d_24_source_34_pat_size_3 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_34_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_34_pat_size_buf_0 <= _source_stream_conv2d_24_source_34_pat_size_0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_34_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_34_pat_size_buf_1 <= _source_stream_conv2d_24_source_34_pat_size_1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_34_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_34_pat_size_buf_2 <= _source_stream_conv2d_24_source_34_pat_size_2;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_34_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_34_pat_size_buf_3 <= _source_stream_conv2d_24_source_34_pat_size_3;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_34_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_34_pat_stride_buf_0 <= _source_stream_conv2d_24_source_34_pat_stride_0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_34_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_34_pat_stride_buf_1 <= _source_stream_conv2d_24_source_34_pat_stride_1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_34_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_34_pat_stride_buf_2 <= _source_stream_conv2d_24_source_34_pat_stride_2;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_34_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_34_pat_stride_buf_3 <= _source_stream_conv2d_24_source_34_pat_stride_3;
      end 
      if(_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_busy && _stream_conv2d_24_is_root) begin
        __variable_wdata_597 <= _stream_conv2d_24_source_34_source_ram_rdata;
      end 
      if((_stream_conv2d_24_source_34_source_pat_fsm_16 == 1) && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_34_idle <= 0;
        _stream_conv2d_24_source_34_source_ram_raddr <= _stream_conv2d_24_source_34_source_pat_all_offset;
        _stream_conv2d_24_source_34_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_24_source_34_source_pat_fsm_16 == 1) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_34_pat_cur_offset_0 <= _source_stream_conv2d_24_source_34_pat_cur_offset_0 + _source_stream_conv2d_24_source_34_pat_stride_buf_0;
        _source_stream_conv2d_24_source_34_pat_count_0 <= _source_stream_conv2d_24_source_34_pat_count_0 - 1;
      end 
      if((_stream_conv2d_24_source_34_source_pat_fsm_16 == 1) && (_source_stream_conv2d_24_source_34_pat_count_0 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_34_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_24_source_34_pat_count_0 <= _source_stream_conv2d_24_source_34_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_24_source_34_source_pat_fsm_16 == 1) && (_source_stream_conv2d_24_source_34_pat_count_0 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_34_pat_cur_offset_1 <= _source_stream_conv2d_24_source_34_pat_cur_offset_1 + _source_stream_conv2d_24_source_34_pat_stride_buf_1;
        _source_stream_conv2d_24_source_34_pat_count_1 <= _source_stream_conv2d_24_source_34_pat_count_1 - 1;
      end 
      if((_stream_conv2d_24_source_34_source_pat_fsm_16 == 1) && (_source_stream_conv2d_24_source_34_pat_count_0 == 0) && (_source_stream_conv2d_24_source_34_pat_count_1 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_34_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_24_source_34_pat_count_1 <= _source_stream_conv2d_24_source_34_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_24_source_34_source_pat_fsm_16 == 1) && ((_source_stream_conv2d_24_source_34_pat_count_0 == 0) && (_source_stream_conv2d_24_source_34_pat_count_1 == 0)) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_34_pat_cur_offset_2 <= _source_stream_conv2d_24_source_34_pat_cur_offset_2 + _source_stream_conv2d_24_source_34_pat_stride_buf_2;
        _source_stream_conv2d_24_source_34_pat_count_2 <= _source_stream_conv2d_24_source_34_pat_count_2 - 1;
      end 
      if((_stream_conv2d_24_source_34_source_pat_fsm_16 == 1) && ((_source_stream_conv2d_24_source_34_pat_count_0 == 0) && (_source_stream_conv2d_24_source_34_pat_count_1 == 0)) && (_source_stream_conv2d_24_source_34_pat_count_2 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_34_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_24_source_34_pat_count_2 <= _source_stream_conv2d_24_source_34_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_24_source_34_source_pat_fsm_16 == 1) && ((_source_stream_conv2d_24_source_34_pat_count_0 == 0) && (_source_stream_conv2d_24_source_34_pat_count_1 == 0) && (_source_stream_conv2d_24_source_34_pat_count_2 == 0)) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_34_pat_cur_offset_3 <= _source_stream_conv2d_24_source_34_pat_cur_offset_3 + _source_stream_conv2d_24_source_34_pat_stride_buf_3;
        _source_stream_conv2d_24_source_34_pat_count_3 <= _source_stream_conv2d_24_source_34_pat_count_3 - 1;
      end 
      if((_stream_conv2d_24_source_34_source_pat_fsm_16 == 1) && ((_source_stream_conv2d_24_source_34_pat_count_0 == 0) && (_source_stream_conv2d_24_source_34_pat_count_1 == 0) && (_source_stream_conv2d_24_source_34_pat_count_2 == 0)) && (_source_stream_conv2d_24_source_34_pat_count_3 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_34_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_24_source_34_pat_count_3 <= _source_stream_conv2d_24_source_34_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_24_source_34_source_pat_fsm_16 == 1) && _stream_conv2d_24_source_stop && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_34_source_ram_renable <= 0;
        _stream_conv2d_24_source_34_idle <= 1;
      end 
      if((_stream_conv2d_24_source_34_source_pat_fsm_16 == 2) && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_34_source_ram_renable <= 0;
        _stream_conv2d_24_source_34_idle <= 1;
      end 
      if(_set_flag_625) begin
        _stream_conv2d_24_source_35_source_mode <= 5'b10;
        _stream_conv2d_24_source_35_source_offset <= conv2d_24_filter_page_comp_offset_buf;
      end 
      if(_set_flag_625) begin
        _source_stream_conv2d_24_source_35_pat_size_0 <= cparam_conv2d_24_stream_reduce_size;
        _source_stream_conv2d_24_source_35_pat_stride_0 <= 1;
      end 
      if(_set_flag_625) begin
        _source_stream_conv2d_24_source_35_pat_size_1 <= conv2d_24_next_stream_num_ops;
        _source_stream_conv2d_24_source_35_pat_stride_1 <= cparam_conv2d_24_stream_aligned_reduce_size;
      end 
      if(_set_flag_625) begin
        _source_stream_conv2d_24_source_35_pat_size_2 <= 1;
        _source_stream_conv2d_24_source_35_pat_stride_2 <= 0;
      end 
      if(_set_flag_625) begin
        _source_stream_conv2d_24_source_35_pat_size_3 <= 1;
        _source_stream_conv2d_24_source_35_pat_stride_3 <= 0;
      end 
      if(_set_flag_625) begin
        _stream_conv2d_24_source_35_source_sel <= 18;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_35_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_35_source_offset_buf <= _stream_conv2d_24_source_35_source_offset;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_35_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_35_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_35_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_35_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_35_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_35_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_35_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_35_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_35_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_35_pat_count_0 <= _source_stream_conv2d_24_source_35_pat_size_0 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_35_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_35_pat_count_1 <= _source_stream_conv2d_24_source_35_pat_size_1 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_35_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_35_pat_count_2 <= _source_stream_conv2d_24_source_35_pat_size_2 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_35_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_35_pat_count_3 <= _source_stream_conv2d_24_source_35_pat_size_3 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_35_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_35_pat_size_buf_0 <= _source_stream_conv2d_24_source_35_pat_size_0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_35_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_35_pat_size_buf_1 <= _source_stream_conv2d_24_source_35_pat_size_1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_35_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_35_pat_size_buf_2 <= _source_stream_conv2d_24_source_35_pat_size_2;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_35_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_35_pat_size_buf_3 <= _source_stream_conv2d_24_source_35_pat_size_3;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_35_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_35_pat_stride_buf_0 <= _source_stream_conv2d_24_source_35_pat_stride_0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_35_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_35_pat_stride_buf_1 <= _source_stream_conv2d_24_source_35_pat_stride_1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_35_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_35_pat_stride_buf_2 <= _source_stream_conv2d_24_source_35_pat_stride_2;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_35_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_35_pat_stride_buf_3 <= _source_stream_conv2d_24_source_35_pat_stride_3;
      end 
      if(_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_busy && _stream_conv2d_24_is_root) begin
        __variable_wdata_598 <= _stream_conv2d_24_source_35_source_ram_rdata;
      end 
      if((_stream_conv2d_24_source_35_source_pat_fsm_17 == 1) && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_35_idle <= 0;
        _stream_conv2d_24_source_35_source_ram_raddr <= _stream_conv2d_24_source_35_source_pat_all_offset;
        _stream_conv2d_24_source_35_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_24_source_35_source_pat_fsm_17 == 1) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_35_pat_cur_offset_0 <= _source_stream_conv2d_24_source_35_pat_cur_offset_0 + _source_stream_conv2d_24_source_35_pat_stride_buf_0;
        _source_stream_conv2d_24_source_35_pat_count_0 <= _source_stream_conv2d_24_source_35_pat_count_0 - 1;
      end 
      if((_stream_conv2d_24_source_35_source_pat_fsm_17 == 1) && (_source_stream_conv2d_24_source_35_pat_count_0 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_35_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_24_source_35_pat_count_0 <= _source_stream_conv2d_24_source_35_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_24_source_35_source_pat_fsm_17 == 1) && (_source_stream_conv2d_24_source_35_pat_count_0 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_35_pat_cur_offset_1 <= _source_stream_conv2d_24_source_35_pat_cur_offset_1 + _source_stream_conv2d_24_source_35_pat_stride_buf_1;
        _source_stream_conv2d_24_source_35_pat_count_1 <= _source_stream_conv2d_24_source_35_pat_count_1 - 1;
      end 
      if((_stream_conv2d_24_source_35_source_pat_fsm_17 == 1) && (_source_stream_conv2d_24_source_35_pat_count_0 == 0) && (_source_stream_conv2d_24_source_35_pat_count_1 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_35_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_24_source_35_pat_count_1 <= _source_stream_conv2d_24_source_35_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_24_source_35_source_pat_fsm_17 == 1) && ((_source_stream_conv2d_24_source_35_pat_count_0 == 0) && (_source_stream_conv2d_24_source_35_pat_count_1 == 0)) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_35_pat_cur_offset_2 <= _source_stream_conv2d_24_source_35_pat_cur_offset_2 + _source_stream_conv2d_24_source_35_pat_stride_buf_2;
        _source_stream_conv2d_24_source_35_pat_count_2 <= _source_stream_conv2d_24_source_35_pat_count_2 - 1;
      end 
      if((_stream_conv2d_24_source_35_source_pat_fsm_17 == 1) && ((_source_stream_conv2d_24_source_35_pat_count_0 == 0) && (_source_stream_conv2d_24_source_35_pat_count_1 == 0)) && (_source_stream_conv2d_24_source_35_pat_count_2 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_35_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_24_source_35_pat_count_2 <= _source_stream_conv2d_24_source_35_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_24_source_35_source_pat_fsm_17 == 1) && ((_source_stream_conv2d_24_source_35_pat_count_0 == 0) && (_source_stream_conv2d_24_source_35_pat_count_1 == 0) && (_source_stream_conv2d_24_source_35_pat_count_2 == 0)) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_35_pat_cur_offset_3 <= _source_stream_conv2d_24_source_35_pat_cur_offset_3 + _source_stream_conv2d_24_source_35_pat_stride_buf_3;
        _source_stream_conv2d_24_source_35_pat_count_3 <= _source_stream_conv2d_24_source_35_pat_count_3 - 1;
      end 
      if((_stream_conv2d_24_source_35_source_pat_fsm_17 == 1) && ((_source_stream_conv2d_24_source_35_pat_count_0 == 0) && (_source_stream_conv2d_24_source_35_pat_count_1 == 0) && (_source_stream_conv2d_24_source_35_pat_count_2 == 0)) && (_source_stream_conv2d_24_source_35_pat_count_3 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_35_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_24_source_35_pat_count_3 <= _source_stream_conv2d_24_source_35_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_24_source_35_source_pat_fsm_17 == 1) && _stream_conv2d_24_source_stop && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_35_source_ram_renable <= 0;
        _stream_conv2d_24_source_35_idle <= 1;
      end 
      if((_stream_conv2d_24_source_35_source_pat_fsm_17 == 2) && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_35_source_ram_renable <= 0;
        _stream_conv2d_24_source_35_idle <= 1;
      end 
      if(_set_flag_638) begin
        _stream_conv2d_24_source_36_source_mode <= 5'b10;
        _stream_conv2d_24_source_36_source_offset <= conv2d_24_filter_page_comp_offset_buf;
      end 
      if(_set_flag_638) begin
        _source_stream_conv2d_24_source_36_pat_size_0 <= cparam_conv2d_24_stream_reduce_size;
        _source_stream_conv2d_24_source_36_pat_stride_0 <= 1;
      end 
      if(_set_flag_638) begin
        _source_stream_conv2d_24_source_36_pat_size_1 <= conv2d_24_next_stream_num_ops;
        _source_stream_conv2d_24_source_36_pat_stride_1 <= cparam_conv2d_24_stream_aligned_reduce_size;
      end 
      if(_set_flag_638) begin
        _source_stream_conv2d_24_source_36_pat_size_2 <= 1;
        _source_stream_conv2d_24_source_36_pat_stride_2 <= 0;
      end 
      if(_set_flag_638) begin
        _source_stream_conv2d_24_source_36_pat_size_3 <= 1;
        _source_stream_conv2d_24_source_36_pat_stride_3 <= 0;
      end 
      if(_set_flag_638) begin
        _stream_conv2d_24_source_36_source_sel <= 19;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_36_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_36_source_offset_buf <= _stream_conv2d_24_source_36_source_offset;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_36_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_36_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_36_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_36_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_36_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_36_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_36_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_36_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_36_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_36_pat_count_0 <= _source_stream_conv2d_24_source_36_pat_size_0 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_36_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_36_pat_count_1 <= _source_stream_conv2d_24_source_36_pat_size_1 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_36_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_36_pat_count_2 <= _source_stream_conv2d_24_source_36_pat_size_2 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_36_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_36_pat_count_3 <= _source_stream_conv2d_24_source_36_pat_size_3 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_36_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_36_pat_size_buf_0 <= _source_stream_conv2d_24_source_36_pat_size_0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_36_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_36_pat_size_buf_1 <= _source_stream_conv2d_24_source_36_pat_size_1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_36_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_36_pat_size_buf_2 <= _source_stream_conv2d_24_source_36_pat_size_2;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_36_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_36_pat_size_buf_3 <= _source_stream_conv2d_24_source_36_pat_size_3;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_36_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_36_pat_stride_buf_0 <= _source_stream_conv2d_24_source_36_pat_stride_0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_36_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_36_pat_stride_buf_1 <= _source_stream_conv2d_24_source_36_pat_stride_1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_36_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_36_pat_stride_buf_2 <= _source_stream_conv2d_24_source_36_pat_stride_2;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_36_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_36_pat_stride_buf_3 <= _source_stream_conv2d_24_source_36_pat_stride_3;
      end 
      if(_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_busy && _stream_conv2d_24_is_root) begin
        __variable_wdata_599 <= _stream_conv2d_24_source_36_source_ram_rdata;
      end 
      if((_stream_conv2d_24_source_36_source_pat_fsm_18 == 1) && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_36_idle <= 0;
        _stream_conv2d_24_source_36_source_ram_raddr <= _stream_conv2d_24_source_36_source_pat_all_offset;
        _stream_conv2d_24_source_36_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_24_source_36_source_pat_fsm_18 == 1) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_36_pat_cur_offset_0 <= _source_stream_conv2d_24_source_36_pat_cur_offset_0 + _source_stream_conv2d_24_source_36_pat_stride_buf_0;
        _source_stream_conv2d_24_source_36_pat_count_0 <= _source_stream_conv2d_24_source_36_pat_count_0 - 1;
      end 
      if((_stream_conv2d_24_source_36_source_pat_fsm_18 == 1) && (_source_stream_conv2d_24_source_36_pat_count_0 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_36_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_24_source_36_pat_count_0 <= _source_stream_conv2d_24_source_36_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_24_source_36_source_pat_fsm_18 == 1) && (_source_stream_conv2d_24_source_36_pat_count_0 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_36_pat_cur_offset_1 <= _source_stream_conv2d_24_source_36_pat_cur_offset_1 + _source_stream_conv2d_24_source_36_pat_stride_buf_1;
        _source_stream_conv2d_24_source_36_pat_count_1 <= _source_stream_conv2d_24_source_36_pat_count_1 - 1;
      end 
      if((_stream_conv2d_24_source_36_source_pat_fsm_18 == 1) && (_source_stream_conv2d_24_source_36_pat_count_0 == 0) && (_source_stream_conv2d_24_source_36_pat_count_1 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_36_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_24_source_36_pat_count_1 <= _source_stream_conv2d_24_source_36_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_24_source_36_source_pat_fsm_18 == 1) && ((_source_stream_conv2d_24_source_36_pat_count_0 == 0) && (_source_stream_conv2d_24_source_36_pat_count_1 == 0)) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_36_pat_cur_offset_2 <= _source_stream_conv2d_24_source_36_pat_cur_offset_2 + _source_stream_conv2d_24_source_36_pat_stride_buf_2;
        _source_stream_conv2d_24_source_36_pat_count_2 <= _source_stream_conv2d_24_source_36_pat_count_2 - 1;
      end 
      if((_stream_conv2d_24_source_36_source_pat_fsm_18 == 1) && ((_source_stream_conv2d_24_source_36_pat_count_0 == 0) && (_source_stream_conv2d_24_source_36_pat_count_1 == 0)) && (_source_stream_conv2d_24_source_36_pat_count_2 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_36_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_24_source_36_pat_count_2 <= _source_stream_conv2d_24_source_36_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_24_source_36_source_pat_fsm_18 == 1) && ((_source_stream_conv2d_24_source_36_pat_count_0 == 0) && (_source_stream_conv2d_24_source_36_pat_count_1 == 0) && (_source_stream_conv2d_24_source_36_pat_count_2 == 0)) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_36_pat_cur_offset_3 <= _source_stream_conv2d_24_source_36_pat_cur_offset_3 + _source_stream_conv2d_24_source_36_pat_stride_buf_3;
        _source_stream_conv2d_24_source_36_pat_count_3 <= _source_stream_conv2d_24_source_36_pat_count_3 - 1;
      end 
      if((_stream_conv2d_24_source_36_source_pat_fsm_18 == 1) && ((_source_stream_conv2d_24_source_36_pat_count_0 == 0) && (_source_stream_conv2d_24_source_36_pat_count_1 == 0) && (_source_stream_conv2d_24_source_36_pat_count_2 == 0)) && (_source_stream_conv2d_24_source_36_pat_count_3 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_36_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_24_source_36_pat_count_3 <= _source_stream_conv2d_24_source_36_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_24_source_36_source_pat_fsm_18 == 1) && _stream_conv2d_24_source_stop && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_36_source_ram_renable <= 0;
        _stream_conv2d_24_source_36_idle <= 1;
      end 
      if((_stream_conv2d_24_source_36_source_pat_fsm_18 == 2) && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_36_source_ram_renable <= 0;
        _stream_conv2d_24_source_36_idle <= 1;
      end 
      if(_set_flag_651) begin
        _stream_conv2d_24_source_37_source_mode <= 5'b10;
        _stream_conv2d_24_source_37_source_offset <= conv2d_24_filter_page_comp_offset_buf;
      end 
      if(_set_flag_651) begin
        _source_stream_conv2d_24_source_37_pat_size_0 <= cparam_conv2d_24_stream_reduce_size;
        _source_stream_conv2d_24_source_37_pat_stride_0 <= 1;
      end 
      if(_set_flag_651) begin
        _source_stream_conv2d_24_source_37_pat_size_1 <= conv2d_24_next_stream_num_ops;
        _source_stream_conv2d_24_source_37_pat_stride_1 <= cparam_conv2d_24_stream_aligned_reduce_size;
      end 
      if(_set_flag_651) begin
        _source_stream_conv2d_24_source_37_pat_size_2 <= 1;
        _source_stream_conv2d_24_source_37_pat_stride_2 <= 0;
      end 
      if(_set_flag_651) begin
        _source_stream_conv2d_24_source_37_pat_size_3 <= 1;
        _source_stream_conv2d_24_source_37_pat_stride_3 <= 0;
      end 
      if(_set_flag_651) begin
        _stream_conv2d_24_source_37_source_sel <= 20;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_37_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_37_source_offset_buf <= _stream_conv2d_24_source_37_source_offset;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_37_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_37_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_37_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_37_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_37_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_37_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_37_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_37_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_37_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_37_pat_count_0 <= _source_stream_conv2d_24_source_37_pat_size_0 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_37_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_37_pat_count_1 <= _source_stream_conv2d_24_source_37_pat_size_1 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_37_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_37_pat_count_2 <= _source_stream_conv2d_24_source_37_pat_size_2 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_37_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_37_pat_count_3 <= _source_stream_conv2d_24_source_37_pat_size_3 - 1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_37_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_37_pat_size_buf_0 <= _source_stream_conv2d_24_source_37_pat_size_0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_37_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_37_pat_size_buf_1 <= _source_stream_conv2d_24_source_37_pat_size_1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_37_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_37_pat_size_buf_2 <= _source_stream_conv2d_24_source_37_pat_size_2;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_37_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_37_pat_size_buf_3 <= _source_stream_conv2d_24_source_37_pat_size_3;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_37_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_37_pat_stride_buf_0 <= _source_stream_conv2d_24_source_37_pat_stride_0;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_37_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_37_pat_stride_buf_1 <= _source_stream_conv2d_24_source_37_pat_stride_1;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_37_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_37_pat_stride_buf_2 <= _source_stream_conv2d_24_source_37_pat_stride_2;
      end 
      if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_37_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_37_pat_stride_buf_3 <= _source_stream_conv2d_24_source_37_pat_stride_3;
      end 
      if(_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_busy && _stream_conv2d_24_is_root) begin
        __variable_wdata_600 <= _stream_conv2d_24_source_37_source_ram_rdata;
      end 
      if((_stream_conv2d_24_source_37_source_pat_fsm_19 == 1) && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_37_idle <= 0;
        _stream_conv2d_24_source_37_source_ram_raddr <= _stream_conv2d_24_source_37_source_pat_all_offset;
        _stream_conv2d_24_source_37_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_24_source_37_source_pat_fsm_19 == 1) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_37_pat_cur_offset_0 <= _source_stream_conv2d_24_source_37_pat_cur_offset_0 + _source_stream_conv2d_24_source_37_pat_stride_buf_0;
        _source_stream_conv2d_24_source_37_pat_count_0 <= _source_stream_conv2d_24_source_37_pat_count_0 - 1;
      end 
      if((_stream_conv2d_24_source_37_source_pat_fsm_19 == 1) && (_source_stream_conv2d_24_source_37_pat_count_0 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_37_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_24_source_37_pat_count_0 <= _source_stream_conv2d_24_source_37_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_24_source_37_source_pat_fsm_19 == 1) && (_source_stream_conv2d_24_source_37_pat_count_0 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_37_pat_cur_offset_1 <= _source_stream_conv2d_24_source_37_pat_cur_offset_1 + _source_stream_conv2d_24_source_37_pat_stride_buf_1;
        _source_stream_conv2d_24_source_37_pat_count_1 <= _source_stream_conv2d_24_source_37_pat_count_1 - 1;
      end 
      if((_stream_conv2d_24_source_37_source_pat_fsm_19 == 1) && (_source_stream_conv2d_24_source_37_pat_count_0 == 0) && (_source_stream_conv2d_24_source_37_pat_count_1 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_37_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_24_source_37_pat_count_1 <= _source_stream_conv2d_24_source_37_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_24_source_37_source_pat_fsm_19 == 1) && ((_source_stream_conv2d_24_source_37_pat_count_0 == 0) && (_source_stream_conv2d_24_source_37_pat_count_1 == 0)) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_37_pat_cur_offset_2 <= _source_stream_conv2d_24_source_37_pat_cur_offset_2 + _source_stream_conv2d_24_source_37_pat_stride_buf_2;
        _source_stream_conv2d_24_source_37_pat_count_2 <= _source_stream_conv2d_24_source_37_pat_count_2 - 1;
      end 
      if((_stream_conv2d_24_source_37_source_pat_fsm_19 == 1) && ((_source_stream_conv2d_24_source_37_pat_count_0 == 0) && (_source_stream_conv2d_24_source_37_pat_count_1 == 0)) && (_source_stream_conv2d_24_source_37_pat_count_2 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_37_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_24_source_37_pat_count_2 <= _source_stream_conv2d_24_source_37_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_24_source_37_source_pat_fsm_19 == 1) && ((_source_stream_conv2d_24_source_37_pat_count_0 == 0) && (_source_stream_conv2d_24_source_37_pat_count_1 == 0) && (_source_stream_conv2d_24_source_37_pat_count_2 == 0)) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_37_pat_cur_offset_3 <= _source_stream_conv2d_24_source_37_pat_cur_offset_3 + _source_stream_conv2d_24_source_37_pat_stride_buf_3;
        _source_stream_conv2d_24_source_37_pat_count_3 <= _source_stream_conv2d_24_source_37_pat_count_3 - 1;
      end 
      if((_stream_conv2d_24_source_37_source_pat_fsm_19 == 1) && ((_source_stream_conv2d_24_source_37_pat_count_0 == 0) && (_source_stream_conv2d_24_source_37_pat_count_1 == 0) && (_source_stream_conv2d_24_source_37_pat_count_2 == 0)) && (_source_stream_conv2d_24_source_37_pat_count_3 == 0) && _stream_conv2d_24_stream_oready) begin
        _source_stream_conv2d_24_source_37_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_24_source_37_pat_count_3 <= _source_stream_conv2d_24_source_37_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_24_source_37_source_pat_fsm_19 == 1) && _stream_conv2d_24_source_stop && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_37_source_ram_renable <= 0;
        _stream_conv2d_24_source_37_idle <= 1;
      end 
      if((_stream_conv2d_24_source_37_source_pat_fsm_19 == 2) && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_source_37_source_ram_renable <= 0;
        _stream_conv2d_24_source_37_idle <= 1;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_665 <= _set_flag_664;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_666 <= _tmp_665;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_667 <= _tmp_666;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_668 <= _tmp_667;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_669 <= _tmp_668;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_670 <= _tmp_669;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_671 <= _tmp_670;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_672 <= _tmp_671;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_673 <= _tmp_672;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_674 <= _tmp_673;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_675 <= _tmp_674;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_676 <= _tmp_675;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_677 <= _tmp_676;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_678 <= _tmp_677;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_679 <= _tmp_678;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_680 <= _tmp_679;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_681 <= _tmp_680;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_682 <= _tmp_681;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_683 <= _tmp_682;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_684 <= _tmp_683;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_685 <= _tmp_684;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_686 <= _tmp_685;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_687 <= _tmp_686;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_688 <= _tmp_687;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_689 <= _tmp_688;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_690 <= _tmp_689;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_691 <= _tmp_690;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_692 <= _tmp_691;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_693 <= _tmp_692;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_694 <= _tmp_693;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_695 <= _tmp_694;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_696 <= _tmp_695;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_697 <= _tmp_696;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_700 <= _tmp_699;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_701 <= _tmp_700;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_702 <= _tmp_701;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_703 <= _tmp_702;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_704 <= _tmp_703;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_705 <= _tmp_704;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_706 <= _tmp_705;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_707 <= _tmp_706;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_708 <= _tmp_707;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_709 <= _tmp_708;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_710 <= _tmp_709;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_711 <= _tmp_710;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_712 <= _tmp_711;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_713 <= _tmp_712;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_714 <= _tmp_713;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_715 <= _tmp_714;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_716 <= _tmp_715;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_717 <= _tmp_716;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_718 <= _tmp_717;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_719 <= _tmp_718;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_720 <= _tmp_719;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_721 <= _tmp_720;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_722 <= _tmp_721;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_723 <= _tmp_722;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_724 <= _tmp_723;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_725 <= _tmp_724;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_726 <= _tmp_725;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_727 <= _tmp_726;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_728 <= _tmp_727;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_729 <= _tmp_728;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_730 <= _tmp_729;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_731 <= _tmp_730;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_732 <= _tmp_731;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_733 <= conv2d_24_next_stream_num_ops;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_734 <= _tmp_733;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_735 <= _tmp_734;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_736 <= _tmp_735;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_737 <= _tmp_736;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_738 <= _tmp_737;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_739 <= _tmp_738;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_740 <= _tmp_739;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_741 <= _tmp_740;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_742 <= _tmp_741;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_743 <= _tmp_742;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_744 <= _tmp_743;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_745 <= _tmp_744;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_746 <= _tmp_745;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_747 <= _tmp_746;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_748 <= _tmp_747;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_749 <= _tmp_748;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_750 <= _tmp_749;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_751 <= _tmp_750;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_752 <= _tmp_751;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_753 <= _tmp_752;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_754 <= _tmp_753;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_755 <= _tmp_754;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_756 <= _tmp_755;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_757 <= _tmp_756;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_758 <= _tmp_757;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_759 <= _tmp_758;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_760 <= _tmp_759;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_761 <= _tmp_760;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_762 <= _tmp_761;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_763 <= _tmp_762;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_764 <= _tmp_763;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_765 <= _tmp_764;
      end 
      if(_tmp_697) begin
        _stream_conv2d_24_sink_50_sink_mode <= 5'b1;
        _stream_conv2d_24_sink_50_sink_offset <= _tmp_732;
        _stream_conv2d_24_sink_50_sink_size <= _tmp_765;
        _stream_conv2d_24_sink_50_sink_stride <= 1;
      end 
      if(_tmp_697) begin
        _stream_conv2d_24_sink_50_sink_sel <= 21;
      end 
      if(_stream_conv2d_24_sink_start && _stream_conv2d_24_sink_50_sink_mode & 5'b1 && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_sink_50_sink_offset_buf <= _stream_conv2d_24_sink_50_sink_offset;
        _stream_conv2d_24_sink_50_sink_size_buf <= _stream_conv2d_24_sink_50_sink_size;
        _stream_conv2d_24_sink_50_sink_stride_buf <= _stream_conv2d_24_sink_50_sink_stride;
      end 
      if((_stream_conv2d_24_sink_50_sink_fsm_20 == 1) && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_sink_50_sink_waddr <= _stream_conv2d_24_sink_50_sink_offset_buf - _stream_conv2d_24_sink_50_sink_stride_buf;
        _stream_conv2d_24_sink_50_sink_count <= _stream_conv2d_24_sink_50_sink_size_buf;
      end 
      if((_stream_conv2d_24_sink_50_sink_fsm_20 == 2) && stream_conv2d_24_sink_51_data && _stream_conv2d_24_stream_oready) begin
        _stream_conv2d_24_sink_50_sink_waddr <= _stream_conv2d_24_sink_50_sink_waddr + _stream_conv2d_24_sink_50_sink_stride_buf;
        _stream_conv2d_24_sink_50_sink_wdata <= stream_conv2d_24_sink_50_data;
        _stream_conv2d_24_sink_50_sink_wenable <= 1;
        _stream_conv2d_24_sink_50_sink_count <= _stream_conv2d_24_sink_50_sink_count - 1;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1156 <= _stream_conv2d_24_source_start;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1157 <= _tmp_1156;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1158 <= _tmp_1157;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1159 <= _stream_conv2d_24_source_start;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1160 <= _tmp_1159;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1161 <= _tmp_1160;
      end 
      if(_stream_conv2d_24_stream_oready && _tmp_1161) begin
        __variable_wdata_309 <= 1;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1162 <= _stream_conv2d_24_source_start;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1163 <= _tmp_1162;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1164 <= _tmp_1163;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1165 <= _tmp_1164;
      end 
      if(_stream_conv2d_24_stream_oready && _tmp_1165) begin
        __variable_wdata_309 <= 0;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1168 <= _tmp_1167;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1171 <= _tmp_1170;
      end 
      if(_stream_conv2d_24_stream_oready && _tmp_1171) begin
        __variable_wdata_309 <= 1;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1172 <= _stream_conv2d_24_source_start;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1173 <= _tmp_1172;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1174 <= _tmp_1173;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1175 <= _tmp_1174;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1176 <= _tmp_1175;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1177 <= _tmp_1176;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1178 <= _tmp_1177;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1179 <= _tmp_1178;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1180 <= _tmp_1179;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1181 <= _tmp_1180;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1182 <= _tmp_1181;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1183 <= _tmp_1182;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1184 <= _tmp_1183;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1185 <= _tmp_1184;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1186 <= _tmp_1185;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1187 <= _tmp_1186;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1188 <= _tmp_1187;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1189 <= _tmp_1188;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1190 <= _tmp_1189;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1191 <= _tmp_1190;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1192 <= _tmp_1191;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1193 <= _tmp_1192;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1194 <= _tmp_1193;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1195 <= _tmp_1194;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1196 <= _tmp_1195;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1197 <= _tmp_1196;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1198 <= _tmp_1197;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1199 <= _tmp_1198;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1200 <= _tmp_1199;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1201 <= _tmp_1200;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1202 <= _tmp_1201;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1203 <= _tmp_1202;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1204 <= _tmp_1203;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1205 <= _stream_conv2d_24_source_stop;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1206 <= _tmp_1205;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1207 <= _tmp_1206;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1208 <= _tmp_1207;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1209 <= _tmp_1208;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1210 <= _tmp_1209;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1211 <= _tmp_1210;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1212 <= _tmp_1211;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1213 <= _tmp_1212;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1214 <= _tmp_1213;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1215 <= _tmp_1214;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1216 <= _tmp_1215;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1217 <= _tmp_1216;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1218 <= _tmp_1217;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1219 <= _tmp_1218;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1220 <= _tmp_1219;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1221 <= _tmp_1220;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1222 <= _tmp_1221;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1223 <= _tmp_1222;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1224 <= _tmp_1223;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1225 <= _tmp_1224;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1226 <= _tmp_1225;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1227 <= _tmp_1226;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1228 <= _tmp_1227;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1229 <= _tmp_1228;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1230 <= _tmp_1229;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1231 <= _tmp_1230;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1232 <= _tmp_1231;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1233 <= _tmp_1232;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1234 <= _tmp_1233;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1235 <= _tmp_1234;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1236 <= _tmp_1235;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1237 <= _tmp_1236;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1238 <= _stream_conv2d_24_source_busy;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1239 <= _tmp_1238;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1240 <= _tmp_1239;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1241 <= _tmp_1240;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1242 <= _tmp_1241;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1243 <= _tmp_1242;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1244 <= _tmp_1243;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1245 <= _tmp_1244;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1246 <= _tmp_1245;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1247 <= _tmp_1246;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1248 <= _tmp_1247;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1249 <= _tmp_1248;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1250 <= _tmp_1249;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1251 <= _tmp_1250;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1252 <= _tmp_1251;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1253 <= _tmp_1252;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1254 <= _tmp_1253;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1255 <= _tmp_1254;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1256 <= _tmp_1255;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1257 <= _tmp_1256;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1258 <= _tmp_1257;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1259 <= _tmp_1258;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1260 <= _tmp_1259;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1261 <= _tmp_1260;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1262 <= _tmp_1261;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1263 <= _tmp_1262;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1264 <= _tmp_1263;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1265 <= _tmp_1264;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1266 <= _tmp_1265;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1267 <= _tmp_1266;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1268 <= _tmp_1267;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1269 <= _tmp_1268;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1270 <= _tmp_1269;
      end 
      if(_stream_conv2d_24_stream_oready) begin
        _tmp_1271 <= _stream_conv2d_24_sink_busy;
      end 
      if(!_stream_conv2d_24_sink_busy && _tmp_1271) begin
        _stream_conv2d_24_busy_reg <= 0;
      end 
      if(_stream_conv2d_24_source_busy) begin
        _stream_conv2d_24_busy_reg <= 1;
      end 
    end
  end

  localparam _stream_conv2d_24_fsm_1 = 1;
  localparam _stream_conv2d_24_fsm_2 = 2;
  localparam _stream_conv2d_24_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_24_fsm <= _stream_conv2d_24_fsm_init;
      _stream_conv2d_24_source_start <= 0;
      _stream_conv2d_24_source_busy <= 0;
      _stream_conv2d_24_stream_ivalid <= 0;
    end else begin
      if(_stream_conv2d_24_stream_oready && _tmp_1158) begin
        _stream_conv2d_24_stream_ivalid <= 1;
      end 
      if(_stream_conv2d_24_stream_oready && _tmp_1168) begin
        _stream_conv2d_24_stream_ivalid <= 0;
      end 
      case(_stream_conv2d_24_fsm)
        _stream_conv2d_24_fsm_init: begin
          if(_stream_conv2d_24_run_flag) begin
            _stream_conv2d_24_source_start <= 1;
          end 
          if(_stream_conv2d_24_run_flag) begin
            _stream_conv2d_24_fsm <= _stream_conv2d_24_fsm_1;
          end 
        end
        _stream_conv2d_24_fsm_1: begin
          if(_stream_conv2d_24_source_start && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_start <= 0;
            _stream_conv2d_24_source_busy <= 1;
          end 
          if(_stream_conv2d_24_source_start && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_fsm <= _stream_conv2d_24_fsm_2;
          end 
        end
        _stream_conv2d_24_fsm_2: begin
          if(_stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_fsm <= _stream_conv2d_24_fsm_3;
          end 
        end
        _stream_conv2d_24_fsm_3: begin
          if(_stream_conv2d_24_stream_oready && (_stream_conv2d_24_source_11_idle && _stream_conv2d_24_source_13_idle && _stream_conv2d_24_source_15_idle && _stream_conv2d_24_source_20_idle && _stream_conv2d_24_source_21_idle && _stream_conv2d_24_source_22_idle && _stream_conv2d_24_source_23_idle && _stream_conv2d_24_source_24_idle && _stream_conv2d_24_source_25_idle && _stream_conv2d_24_source_26_idle && _stream_conv2d_24_source_27_idle && _stream_conv2d_24_source_28_idle && _stream_conv2d_24_source_29_idle && _stream_conv2d_24_source_30_idle && _stream_conv2d_24_source_31_idle && _stream_conv2d_24_source_32_idle && _stream_conv2d_24_source_33_idle && _stream_conv2d_24_source_34_idle && _stream_conv2d_24_source_35_idle && _stream_conv2d_24_source_36_idle && _stream_conv2d_24_source_37_idle && _stream_conv2d_24_source_7_idle && _stream_conv2d_24_source_9_idle && (_stream_conv2d_24_fsm == 3))) begin
            _stream_conv2d_24_source_busy <= 0;
          end 
          if(_stream_conv2d_24_stream_oready && (_stream_conv2d_24_source_11_idle && _stream_conv2d_24_source_13_idle && _stream_conv2d_24_source_15_idle && _stream_conv2d_24_source_20_idle && _stream_conv2d_24_source_21_idle && _stream_conv2d_24_source_22_idle && _stream_conv2d_24_source_23_idle && _stream_conv2d_24_source_24_idle && _stream_conv2d_24_source_25_idle && _stream_conv2d_24_source_26_idle && _stream_conv2d_24_source_27_idle && _stream_conv2d_24_source_28_idle && _stream_conv2d_24_source_29_idle && _stream_conv2d_24_source_30_idle && _stream_conv2d_24_source_31_idle && _stream_conv2d_24_source_32_idle && _stream_conv2d_24_source_33_idle && _stream_conv2d_24_source_34_idle && _stream_conv2d_24_source_35_idle && _stream_conv2d_24_source_36_idle && _stream_conv2d_24_source_37_idle && _stream_conv2d_24_source_7_idle && _stream_conv2d_24_source_9_idle && (_stream_conv2d_24_fsm == 3)) && _stream_conv2d_24_run_flag) begin
            _stream_conv2d_24_source_start <= 1;
          end 
          if(_stream_conv2d_24_stream_oready && (_stream_conv2d_24_source_11_idle && _stream_conv2d_24_source_13_idle && _stream_conv2d_24_source_15_idle && _stream_conv2d_24_source_20_idle && _stream_conv2d_24_source_21_idle && _stream_conv2d_24_source_22_idle && _stream_conv2d_24_source_23_idle && _stream_conv2d_24_source_24_idle && _stream_conv2d_24_source_25_idle && _stream_conv2d_24_source_26_idle && _stream_conv2d_24_source_27_idle && _stream_conv2d_24_source_28_idle && _stream_conv2d_24_source_29_idle && _stream_conv2d_24_source_30_idle && _stream_conv2d_24_source_31_idle && _stream_conv2d_24_source_32_idle && _stream_conv2d_24_source_33_idle && _stream_conv2d_24_source_34_idle && _stream_conv2d_24_source_35_idle && _stream_conv2d_24_source_36_idle && _stream_conv2d_24_source_37_idle && _stream_conv2d_24_source_7_idle && _stream_conv2d_24_source_9_idle && (_stream_conv2d_24_fsm == 3))) begin
            _stream_conv2d_24_fsm <= _stream_conv2d_24_fsm_init;
          end 
          if(_stream_conv2d_24_stream_oready && (_stream_conv2d_24_source_11_idle && _stream_conv2d_24_source_13_idle && _stream_conv2d_24_source_15_idle && _stream_conv2d_24_source_20_idle && _stream_conv2d_24_source_21_idle && _stream_conv2d_24_source_22_idle && _stream_conv2d_24_source_23_idle && _stream_conv2d_24_source_24_idle && _stream_conv2d_24_source_25_idle && _stream_conv2d_24_source_26_idle && _stream_conv2d_24_source_27_idle && _stream_conv2d_24_source_28_idle && _stream_conv2d_24_source_29_idle && _stream_conv2d_24_source_30_idle && _stream_conv2d_24_source_31_idle && _stream_conv2d_24_source_32_idle && _stream_conv2d_24_source_33_idle && _stream_conv2d_24_source_34_idle && _stream_conv2d_24_source_35_idle && _stream_conv2d_24_source_36_idle && _stream_conv2d_24_source_37_idle && _stream_conv2d_24_source_7_idle && _stream_conv2d_24_source_9_idle && (_stream_conv2d_24_fsm == 3)) && _stream_conv2d_24_run_flag) begin
            _stream_conv2d_24_fsm <= _stream_conv2d_24_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _stream_max_pool_serial_26_source_1_source_ram_renable <= 0;
      _stream_max_pool_serial_26_source_1_source_fifo_deq <= 0;
      _stream_max_pool_serial_26_source_1_idle <= 1;
      _stream_max_pool_serial_26_sink_5_sink_wenable <= 0;
      _stream_max_pool_serial_26_sink_5_sink_fifo_enq <= 0;
      _stream_max_pool_serial_26_sink_6_sink_wenable <= 0;
      _stream_max_pool_serial_26_sink_6_sink_fifo_enq <= 0;
      __stream_max_pool_serial_26_stream_ivalid_1 <= 0;
      __stream_max_pool_serial_26_stream_ivalid_2 <= 0;
      __stream_max_pool_serial_26_stream_ivalid_3 <= 0;
      __stream_max_pool_serial_26_stream_ivalid_4 <= 0;
      __stream_max_pool_serial_26_stream_ivalid_5 <= 0;
      _counter_data_897 <= 1'sd0;
      _counter_count_897 <= 1'sd0;
      __delay_data_1174__variable_895 <= 0;
      __delay_data_1175_reinterpretcast_905 <= 0;
      __delay_data_1177__variable_896 <= 0;
      __delay_data_1180__variable_893 <= 0;
      _pointer_data_900 <= 0;
      __delay_data_1176__delay_1175_reinterpretcast_905 <= 0;
      __delay_data_1178__delay_1177__variable_896 <= 0;
      __delay_data_1181__delay_1180__variable_893 <= 0;
      _cond_data_907 <= 0;
      __delay_data_1179__delay_1178__delay_1177__variable_896 <= 0;
      __delay_data_1182__delay_1181__delay_1180__variable_893 <= 0;
      _stream_max_pool_serial_26_parameter_0_next_parameter_data <= 0;
      __variable_wdata_893 <= 0;
      _stream_max_pool_serial_26_parameter_2_next_parameter_data <= 0;
      __variable_wdata_895 <= 0;
      _stream_max_pool_serial_26_source_1_source_mode <= 5'b0;
      _stream_max_pool_serial_26_source_1_source_offset <= 0;
      _source_stream_max_pool_serial_26_source_1_pat_size_0 <= 0;
      _source_stream_max_pool_serial_26_source_1_pat_stride_0 <= 0;
      _source_stream_max_pool_serial_26_source_1_pat_size_1 <= 0;
      _source_stream_max_pool_serial_26_source_1_pat_stride_1 <= 0;
      _source_stream_max_pool_serial_26_source_1_pat_size_2 <= 0;
      _source_stream_max_pool_serial_26_source_1_pat_stride_2 <= 0;
      _source_stream_max_pool_serial_26_source_1_pat_size_3 <= 0;
      _source_stream_max_pool_serial_26_source_1_pat_stride_3 <= 0;
      _stream_max_pool_serial_26_source_1_source_sel <= 0;
      _stream_max_pool_serial_26_source_1_source_offset_buf <= 0;
      _source_stream_max_pool_serial_26_source_1_pat_cur_offset_0 <= 0;
      _source_stream_max_pool_serial_26_source_1_pat_cur_offset_1 <= 0;
      _source_stream_max_pool_serial_26_source_1_pat_cur_offset_2 <= 0;
      _source_stream_max_pool_serial_26_source_1_pat_cur_offset_3 <= 0;
      _source_stream_max_pool_serial_26_source_1_pat_count_0 <= 0;
      _source_stream_max_pool_serial_26_source_1_pat_count_1 <= 0;
      _source_stream_max_pool_serial_26_source_1_pat_count_2 <= 0;
      _source_stream_max_pool_serial_26_source_1_pat_count_3 <= 0;
      _source_stream_max_pool_serial_26_source_1_pat_size_buf_0 <= 0;
      _source_stream_max_pool_serial_26_source_1_pat_size_buf_1 <= 0;
      _source_stream_max_pool_serial_26_source_1_pat_size_buf_2 <= 0;
      _source_stream_max_pool_serial_26_source_1_pat_size_buf_3 <= 0;
      _source_stream_max_pool_serial_26_source_1_pat_stride_buf_0 <= 0;
      _source_stream_max_pool_serial_26_source_1_pat_stride_buf_1 <= 0;
      _source_stream_max_pool_serial_26_source_1_pat_stride_buf_2 <= 0;
      _source_stream_max_pool_serial_26_source_1_pat_stride_buf_3 <= 0;
      __variable_wdata_894 <= 0;
      _stream_max_pool_serial_26_source_1_source_ram_raddr <= 0;
      _tmp_1365 <= 0;
      _tmp_1366 <= 0;
      _tmp_1367 <= 0;
      _tmp_1368 <= 0;
      _tmp_1369 <= 0;
      _tmp_1370 <= 0;
      _tmp_1371 <= 0;
      _tmp_1374 <= 0;
      _tmp_1375 <= 0;
      _tmp_1376 <= 0;
      _tmp_1377 <= 0;
      _tmp_1378 <= 0;
      _tmp_1379 <= 0;
      _tmp_1380 <= 0;
      _tmp_1381 <= 0;
      _tmp_1382 <= 0;
      _tmp_1383 <= 0;
      _tmp_1384 <= 0;
      _tmp_1385 <= 0;
      _tmp_1386 <= 0;
      _tmp_1387 <= 0;
      _stream_max_pool_serial_26_sink_5_sink_mode <= 5'b0;
      _stream_max_pool_serial_26_sink_5_sink_offset <= 0;
      _stream_max_pool_serial_26_sink_5_sink_size <= 0;
      _stream_max_pool_serial_26_sink_5_sink_stride <= 0;
      _stream_max_pool_serial_26_sink_5_sink_sel <= 0;
      _stream_max_pool_serial_26_sink_5_sink_offset_buf <= 0;
      _stream_max_pool_serial_26_sink_5_sink_size_buf <= 0;
      _stream_max_pool_serial_26_sink_5_sink_stride_buf <= 0;
      _stream_max_pool_serial_26_sink_5_sink_waddr <= 0;
      _stream_max_pool_serial_26_sink_5_sink_count <= 0;
      _stream_max_pool_serial_26_sink_5_sink_wdata <= 0;
      _tmp_1410 <= 0;
      _tmp_1411 <= 0;
      _tmp_1412 <= 0;
      _tmp_1413 <= 0;
      _tmp_1414 <= 0;
      _tmp_1415 <= 0;
      __variable_wdata_896 <= 0;
      _tmp_1416 <= 0;
      _tmp_1417 <= 0;
      _tmp_1418 <= 0;
      _tmp_1419 <= 0;
      _tmp_1422 <= 0;
      _tmp_1425 <= 0;
      _tmp_1426 <= 0;
      _tmp_1427 <= 0;
      _tmp_1428 <= 0;
      _tmp_1429 <= 0;
      _tmp_1430 <= 0;
      _tmp_1431 <= 0;
      _tmp_1432 <= 0;
      _tmp_1433 <= 0;
      _tmp_1434 <= 0;
      _tmp_1435 <= 0;
      _tmp_1436 <= 0;
      _tmp_1437 <= 0;
      _tmp_1438 <= 0;
      _tmp_1439 <= 0;
      _tmp_1440 <= 0;
      _tmp_1441 <= 0;
      _tmp_1442 <= 0;
      _tmp_1443 <= 0;
      _tmp_1444 <= 0;
      _tmp_1445 <= 0;
      _tmp_1446 <= 0;
      _tmp_1447 <= 0;
      _stream_max_pool_serial_26_busy_reg <= 0;
    end else begin
      if(_stream_max_pool_serial_26_stream_oready) begin
        _stream_max_pool_serial_26_source_1_source_ram_renable <= 0;
        _stream_max_pool_serial_26_source_1_source_fifo_deq <= 0;
      end 
      _stream_max_pool_serial_26_source_1_idle <= _stream_max_pool_serial_26_source_1_idle;
      if(_stream_max_pool_serial_26_stream_oready) begin
        _stream_max_pool_serial_26_sink_5_sink_wenable <= 0;
        _stream_max_pool_serial_26_sink_5_sink_fifo_enq <= 0;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _stream_max_pool_serial_26_sink_6_sink_wenable <= 0;
        _stream_max_pool_serial_26_sink_6_sink_fifo_enq <= 0;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        __stream_max_pool_serial_26_stream_ivalid_1 <= _stream_max_pool_serial_26_stream_ivalid;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        __stream_max_pool_serial_26_stream_ivalid_2 <= __stream_max_pool_serial_26_stream_ivalid_1;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        __stream_max_pool_serial_26_stream_ivalid_3 <= __stream_max_pool_serial_26_stream_ivalid_2;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        __stream_max_pool_serial_26_stream_ivalid_4 <= __stream_max_pool_serial_26_stream_ivalid_3;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        __stream_max_pool_serial_26_stream_ivalid_5 <= __stream_max_pool_serial_26_stream_ivalid_4;
      end 
      if(_stream_max_pool_serial_26_stream_ivalid && _stream_max_pool_serial_26_stream_oready && _counter_reset_cond_897) begin
        _counter_data_897 <= 1'sd0;
      end 
      if(_stream_max_pool_serial_26_stream_ivalid && _stream_max_pool_serial_26_stream_oready) begin
        _counter_data_897 <= _counter_current_count_897;
      end 
      if(_stream_max_pool_serial_26_stream_ivalid && _stream_max_pool_serial_26_stream_oready) begin
        _counter_count_897 <= (_counter_current_count_897 >= stream_max_pool_serial_26_parameter_0_data - 2'sd1)? _counter_current_count_897 + 2'sd1 - stream_max_pool_serial_26_parameter_0_data : _counter_current_count_897 + 2'sd1;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        __delay_data_1174__variable_895 <= stream_max_pool_serial_26_parameter_2_data;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        __delay_data_1175_reinterpretcast_905 <= _reinterpretcast_data_905;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        __delay_data_1177__variable_896 <= stream_max_pool_serial_26__reduce_reset_data;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        __delay_data_1180__variable_893 <= stream_max_pool_serial_26_parameter_0_data;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _pointer_data_900 <= __delay_data_1174__variable_895[_counter_data_897];
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        __delay_data_1176__delay_1175_reinterpretcast_905 <= __delay_data_1175_reinterpretcast_905;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        __delay_data_1178__delay_1177__variable_896 <= __delay_data_1177__variable_896;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        __delay_data_1181__delay_1180__variable_893 <= __delay_data_1180__variable_893;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _cond_data_907 <= (_pointer_data_900)? -9'sd128 : __delay_data_1176__delay_1175_reinterpretcast_905;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        __delay_data_1179__delay_1178__delay_1177__variable_896 <= __delay_data_1178__delay_1177__variable_896;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        __delay_data_1182__delay_1181__delay_1180__variable_893 <= __delay_data_1181__delay_1180__variable_893;
      end 
      if(_set_flag_1349) begin
        _stream_max_pool_serial_26_parameter_0_next_parameter_data <= 4;
      end 
      if(_stream_max_pool_serial_26_source_start) begin
        __variable_wdata_893 <= _stream_max_pool_serial_26_parameter_0_next_parameter_data;
      end 
      if(_set_flag_1350) begin
        _stream_max_pool_serial_26_parameter_2_next_parameter_data <= max_pool_serial_26_stream_pad_masks;
      end 
      if(_stream_max_pool_serial_26_source_start) begin
        __variable_wdata_895 <= _stream_max_pool_serial_26_parameter_2_next_parameter_data;
      end 
      if(_set_flag_1351) begin
        _stream_max_pool_serial_26_source_1_source_mode <= 5'b10;
        _stream_max_pool_serial_26_source_1_source_offset <= max_pool_serial_26_stream_act_local + max_pool_serial_26_act_page_comp_offset_buf;
      end 
      if(_set_flag_1351) begin
        _source_stream_max_pool_serial_26_source_1_pat_size_0 <= 2;
        _source_stream_max_pool_serial_26_source_1_pat_stride_0 <= cparam_max_pool_serial_26_act_read_block;
      end 
      if(_set_flag_1351) begin
        _source_stream_max_pool_serial_26_source_1_pat_size_1 <= 2;
        _source_stream_max_pool_serial_26_source_1_pat_stride_1 <= cparam_max_pool_serial_26_act_read_size;
      end 
      if(_set_flag_1351) begin
        _source_stream_max_pool_serial_26_source_1_pat_size_2 <= cparam_max_pool_serial_26_stream_size;
        _source_stream_max_pool_serial_26_source_1_pat_stride_2 <= 1;
      end 
      if(_set_flag_1351) begin
        _source_stream_max_pool_serial_26_source_1_pat_size_3 <= 1;
        _source_stream_max_pool_serial_26_source_1_pat_stride_3 <= 0;
      end 
      if(_set_flag_1351) begin
        _stream_max_pool_serial_26_source_1_source_sel <= 1;
      end 
      if(_stream_max_pool_serial_26_source_start && _stream_max_pool_serial_26_source_1_source_mode & 5'b10 && _stream_max_pool_serial_26_stream_oready) begin
        _stream_max_pool_serial_26_source_1_source_offset_buf <= _stream_max_pool_serial_26_source_1_source_offset;
      end 
      if(_stream_max_pool_serial_26_source_start && _stream_max_pool_serial_26_source_1_source_mode & 5'b10 && _stream_max_pool_serial_26_stream_oready) begin
        _source_stream_max_pool_serial_26_source_1_pat_cur_offset_0 <= 0;
      end 
      if(_stream_max_pool_serial_26_source_start && _stream_max_pool_serial_26_source_1_source_mode & 5'b10 && _stream_max_pool_serial_26_stream_oready) begin
        _source_stream_max_pool_serial_26_source_1_pat_cur_offset_1 <= 0;
      end 
      if(_stream_max_pool_serial_26_source_start && _stream_max_pool_serial_26_source_1_source_mode & 5'b10 && _stream_max_pool_serial_26_stream_oready) begin
        _source_stream_max_pool_serial_26_source_1_pat_cur_offset_2 <= 0;
      end 
      if(_stream_max_pool_serial_26_source_start && _stream_max_pool_serial_26_source_1_source_mode & 5'b10 && _stream_max_pool_serial_26_stream_oready) begin
        _source_stream_max_pool_serial_26_source_1_pat_cur_offset_3 <= 0;
      end 
      if(_stream_max_pool_serial_26_source_start && _stream_max_pool_serial_26_source_1_source_mode & 5'b10 && _stream_max_pool_serial_26_stream_oready) begin
        _source_stream_max_pool_serial_26_source_1_pat_count_0 <= _source_stream_max_pool_serial_26_source_1_pat_size_0 - 1;
      end 
      if(_stream_max_pool_serial_26_source_start && _stream_max_pool_serial_26_source_1_source_mode & 5'b10 && _stream_max_pool_serial_26_stream_oready) begin
        _source_stream_max_pool_serial_26_source_1_pat_count_1 <= _source_stream_max_pool_serial_26_source_1_pat_size_1 - 1;
      end 
      if(_stream_max_pool_serial_26_source_start && _stream_max_pool_serial_26_source_1_source_mode & 5'b10 && _stream_max_pool_serial_26_stream_oready) begin
        _source_stream_max_pool_serial_26_source_1_pat_count_2 <= _source_stream_max_pool_serial_26_source_1_pat_size_2 - 1;
      end 
      if(_stream_max_pool_serial_26_source_start && _stream_max_pool_serial_26_source_1_source_mode & 5'b10 && _stream_max_pool_serial_26_stream_oready) begin
        _source_stream_max_pool_serial_26_source_1_pat_count_3 <= _source_stream_max_pool_serial_26_source_1_pat_size_3 - 1;
      end 
      if(_stream_max_pool_serial_26_source_start && _stream_max_pool_serial_26_source_1_source_mode & 5'b10 && _stream_max_pool_serial_26_stream_oready) begin
        _source_stream_max_pool_serial_26_source_1_pat_size_buf_0 <= _source_stream_max_pool_serial_26_source_1_pat_size_0;
      end 
      if(_stream_max_pool_serial_26_source_start && _stream_max_pool_serial_26_source_1_source_mode & 5'b10 && _stream_max_pool_serial_26_stream_oready) begin
        _source_stream_max_pool_serial_26_source_1_pat_size_buf_1 <= _source_stream_max_pool_serial_26_source_1_pat_size_1;
      end 
      if(_stream_max_pool_serial_26_source_start && _stream_max_pool_serial_26_source_1_source_mode & 5'b10 && _stream_max_pool_serial_26_stream_oready) begin
        _source_stream_max_pool_serial_26_source_1_pat_size_buf_2 <= _source_stream_max_pool_serial_26_source_1_pat_size_2;
      end 
      if(_stream_max_pool_serial_26_source_start && _stream_max_pool_serial_26_source_1_source_mode & 5'b10 && _stream_max_pool_serial_26_stream_oready) begin
        _source_stream_max_pool_serial_26_source_1_pat_size_buf_3 <= _source_stream_max_pool_serial_26_source_1_pat_size_3;
      end 
      if(_stream_max_pool_serial_26_source_start && _stream_max_pool_serial_26_source_1_source_mode & 5'b10 && _stream_max_pool_serial_26_stream_oready) begin
        _source_stream_max_pool_serial_26_source_1_pat_stride_buf_0 <= _source_stream_max_pool_serial_26_source_1_pat_stride_0;
      end 
      if(_stream_max_pool_serial_26_source_start && _stream_max_pool_serial_26_source_1_source_mode & 5'b10 && _stream_max_pool_serial_26_stream_oready) begin
        _source_stream_max_pool_serial_26_source_1_pat_stride_buf_1 <= _source_stream_max_pool_serial_26_source_1_pat_stride_1;
      end 
      if(_stream_max_pool_serial_26_source_start && _stream_max_pool_serial_26_source_1_source_mode & 5'b10 && _stream_max_pool_serial_26_stream_oready) begin
        _source_stream_max_pool_serial_26_source_1_pat_stride_buf_2 <= _source_stream_max_pool_serial_26_source_1_pat_stride_2;
      end 
      if(_stream_max_pool_serial_26_source_start && _stream_max_pool_serial_26_source_1_source_mode & 5'b10 && _stream_max_pool_serial_26_stream_oready) begin
        _source_stream_max_pool_serial_26_source_1_pat_stride_buf_3 <= _source_stream_max_pool_serial_26_source_1_pat_stride_3;
      end 
      if(_stream_max_pool_serial_26_stream_oready && _stream_max_pool_serial_26_source_busy && _stream_max_pool_serial_26_is_root) begin
        __variable_wdata_894 <= _stream_max_pool_serial_26_source_1_source_ram_rdata;
      end 
      if((_stream_max_pool_serial_26_source_1_source_pat_fsm_0 == 1) && _stream_max_pool_serial_26_stream_oready) begin
        _stream_max_pool_serial_26_source_1_idle <= 0;
        _stream_max_pool_serial_26_source_1_source_ram_raddr <= _stream_max_pool_serial_26_source_1_source_pat_all_offset;
        _stream_max_pool_serial_26_source_1_source_ram_renable <= 1;
      end 
      if((_stream_max_pool_serial_26_source_1_source_pat_fsm_0 == 1) && _stream_max_pool_serial_26_stream_oready) begin
        _source_stream_max_pool_serial_26_source_1_pat_cur_offset_0 <= _source_stream_max_pool_serial_26_source_1_pat_cur_offset_0 + _source_stream_max_pool_serial_26_source_1_pat_stride_buf_0;
        _source_stream_max_pool_serial_26_source_1_pat_count_0 <= _source_stream_max_pool_serial_26_source_1_pat_count_0 - 1;
      end 
      if((_stream_max_pool_serial_26_source_1_source_pat_fsm_0 == 1) && (_source_stream_max_pool_serial_26_source_1_pat_count_0 == 0) && _stream_max_pool_serial_26_stream_oready) begin
        _source_stream_max_pool_serial_26_source_1_pat_cur_offset_0 <= 0;
        _source_stream_max_pool_serial_26_source_1_pat_count_0 <= _source_stream_max_pool_serial_26_source_1_pat_size_buf_0 - 1;
      end 
      if((_stream_max_pool_serial_26_source_1_source_pat_fsm_0 == 1) && (_source_stream_max_pool_serial_26_source_1_pat_count_0 == 0) && _stream_max_pool_serial_26_stream_oready) begin
        _source_stream_max_pool_serial_26_source_1_pat_cur_offset_1 <= _source_stream_max_pool_serial_26_source_1_pat_cur_offset_1 + _source_stream_max_pool_serial_26_source_1_pat_stride_buf_1;
        _source_stream_max_pool_serial_26_source_1_pat_count_1 <= _source_stream_max_pool_serial_26_source_1_pat_count_1 - 1;
      end 
      if((_stream_max_pool_serial_26_source_1_source_pat_fsm_0 == 1) && (_source_stream_max_pool_serial_26_source_1_pat_count_0 == 0) && (_source_stream_max_pool_serial_26_source_1_pat_count_1 == 0) && _stream_max_pool_serial_26_stream_oready) begin
        _source_stream_max_pool_serial_26_source_1_pat_cur_offset_1 <= 0;
        _source_stream_max_pool_serial_26_source_1_pat_count_1 <= _source_stream_max_pool_serial_26_source_1_pat_size_buf_1 - 1;
      end 
      if((_stream_max_pool_serial_26_source_1_source_pat_fsm_0 == 1) && ((_source_stream_max_pool_serial_26_source_1_pat_count_0 == 0) && (_source_stream_max_pool_serial_26_source_1_pat_count_1 == 0)) && _stream_max_pool_serial_26_stream_oready) begin
        _source_stream_max_pool_serial_26_source_1_pat_cur_offset_2 <= _source_stream_max_pool_serial_26_source_1_pat_cur_offset_2 + _source_stream_max_pool_serial_26_source_1_pat_stride_buf_2;
        _source_stream_max_pool_serial_26_source_1_pat_count_2 <= _source_stream_max_pool_serial_26_source_1_pat_count_2 - 1;
      end 
      if((_stream_max_pool_serial_26_source_1_source_pat_fsm_0 == 1) && ((_source_stream_max_pool_serial_26_source_1_pat_count_0 == 0) && (_source_stream_max_pool_serial_26_source_1_pat_count_1 == 0)) && (_source_stream_max_pool_serial_26_source_1_pat_count_2 == 0) && _stream_max_pool_serial_26_stream_oready) begin
        _source_stream_max_pool_serial_26_source_1_pat_cur_offset_2 <= 0;
        _source_stream_max_pool_serial_26_source_1_pat_count_2 <= _source_stream_max_pool_serial_26_source_1_pat_size_buf_2 - 1;
      end 
      if((_stream_max_pool_serial_26_source_1_source_pat_fsm_0 == 1) && ((_source_stream_max_pool_serial_26_source_1_pat_count_0 == 0) && (_source_stream_max_pool_serial_26_source_1_pat_count_1 == 0) && (_source_stream_max_pool_serial_26_source_1_pat_count_2 == 0)) && _stream_max_pool_serial_26_stream_oready) begin
        _source_stream_max_pool_serial_26_source_1_pat_cur_offset_3 <= _source_stream_max_pool_serial_26_source_1_pat_cur_offset_3 + _source_stream_max_pool_serial_26_source_1_pat_stride_buf_3;
        _source_stream_max_pool_serial_26_source_1_pat_count_3 <= _source_stream_max_pool_serial_26_source_1_pat_count_3 - 1;
      end 
      if((_stream_max_pool_serial_26_source_1_source_pat_fsm_0 == 1) && ((_source_stream_max_pool_serial_26_source_1_pat_count_0 == 0) && (_source_stream_max_pool_serial_26_source_1_pat_count_1 == 0) && (_source_stream_max_pool_serial_26_source_1_pat_count_2 == 0)) && (_source_stream_max_pool_serial_26_source_1_pat_count_3 == 0) && _stream_max_pool_serial_26_stream_oready) begin
        _source_stream_max_pool_serial_26_source_1_pat_cur_offset_3 <= 0;
        _source_stream_max_pool_serial_26_source_1_pat_count_3 <= _source_stream_max_pool_serial_26_source_1_pat_size_buf_3 - 1;
      end 
      if((_stream_max_pool_serial_26_source_1_source_pat_fsm_0 == 1) && _stream_max_pool_serial_26_source_stop && _stream_max_pool_serial_26_stream_oready) begin
        _stream_max_pool_serial_26_source_1_source_ram_renable <= 0;
        _stream_max_pool_serial_26_source_1_idle <= 1;
      end 
      if((_stream_max_pool_serial_26_source_1_source_pat_fsm_0 == 2) && _stream_max_pool_serial_26_stream_oready) begin
        _stream_max_pool_serial_26_source_1_source_ram_renable <= 0;
        _stream_max_pool_serial_26_source_1_idle <= 1;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _tmp_1365 <= _set_flag_1364;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _tmp_1366 <= _tmp_1365;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _tmp_1367 <= _tmp_1366;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _tmp_1368 <= _tmp_1367;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _tmp_1369 <= _tmp_1368;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _tmp_1370 <= _tmp_1369;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _tmp_1371 <= _tmp_1370;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _tmp_1374 <= _tmp_1373;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _tmp_1375 <= _tmp_1374;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _tmp_1376 <= _tmp_1375;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _tmp_1377 <= _tmp_1376;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _tmp_1378 <= _tmp_1377;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _tmp_1379 <= _tmp_1378;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _tmp_1380 <= _tmp_1379;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _tmp_1381 <= cparam_max_pool_serial_26_stream_size;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _tmp_1382 <= _tmp_1381;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _tmp_1383 <= _tmp_1382;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _tmp_1384 <= _tmp_1383;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _tmp_1385 <= _tmp_1384;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _tmp_1386 <= _tmp_1385;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _tmp_1387 <= _tmp_1386;
      end 
      if(_tmp_1371) begin
        _stream_max_pool_serial_26_sink_5_sink_mode <= 5'b1;
        _stream_max_pool_serial_26_sink_5_sink_offset <= _tmp_1380;
        _stream_max_pool_serial_26_sink_5_sink_size <= _tmp_1387;
        _stream_max_pool_serial_26_sink_5_sink_stride <= 1;
      end 
      if(_tmp_1371) begin
        _stream_max_pool_serial_26_sink_5_sink_sel <= 2;
      end 
      if(_stream_max_pool_serial_26_sink_start && _stream_max_pool_serial_26_sink_5_sink_mode & 5'b1 && _stream_max_pool_serial_26_stream_oready) begin
        _stream_max_pool_serial_26_sink_5_sink_offset_buf <= _stream_max_pool_serial_26_sink_5_sink_offset;
        _stream_max_pool_serial_26_sink_5_sink_size_buf <= _stream_max_pool_serial_26_sink_5_sink_size;
        _stream_max_pool_serial_26_sink_5_sink_stride_buf <= _stream_max_pool_serial_26_sink_5_sink_stride;
      end 
      if((_stream_max_pool_serial_26_sink_5_sink_fsm_1 == 1) && _stream_max_pool_serial_26_stream_oready) begin
        _stream_max_pool_serial_26_sink_5_sink_waddr <= _stream_max_pool_serial_26_sink_5_sink_offset_buf - _stream_max_pool_serial_26_sink_5_sink_stride_buf;
        _stream_max_pool_serial_26_sink_5_sink_count <= _stream_max_pool_serial_26_sink_5_sink_size_buf;
      end 
      if((_stream_max_pool_serial_26_sink_5_sink_fsm_1 == 2) && stream_max_pool_serial_26_sink_6_data && _stream_max_pool_serial_26_stream_oready) begin
        _stream_max_pool_serial_26_sink_5_sink_waddr <= _stream_max_pool_serial_26_sink_5_sink_waddr + _stream_max_pool_serial_26_sink_5_sink_stride_buf;
        _stream_max_pool_serial_26_sink_5_sink_wdata <= stream_max_pool_serial_26_sink_5_data;
        _stream_max_pool_serial_26_sink_5_sink_wenable <= 1;
        _stream_max_pool_serial_26_sink_5_sink_count <= _stream_max_pool_serial_26_sink_5_sink_count - 1;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _tmp_1410 <= _stream_max_pool_serial_26_source_start;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _tmp_1411 <= _tmp_1410;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _tmp_1412 <= _tmp_1411;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _tmp_1413 <= _stream_max_pool_serial_26_source_start;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _tmp_1414 <= _tmp_1413;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _tmp_1415 <= _tmp_1414;
      end 
      if(_stream_max_pool_serial_26_stream_oready && _tmp_1415) begin
        __variable_wdata_896 <= 1;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _tmp_1416 <= _stream_max_pool_serial_26_source_start;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _tmp_1417 <= _tmp_1416;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _tmp_1418 <= _tmp_1417;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _tmp_1419 <= _tmp_1418;
      end 
      if(_stream_max_pool_serial_26_stream_oready && _tmp_1419) begin
        __variable_wdata_896 <= 0;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _tmp_1422 <= _tmp_1421;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _tmp_1425 <= _tmp_1424;
      end 
      if(_stream_max_pool_serial_26_stream_oready && _tmp_1425) begin
        __variable_wdata_896 <= 1;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _tmp_1426 <= _stream_max_pool_serial_26_source_start;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _tmp_1427 <= _tmp_1426;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _tmp_1428 <= _tmp_1427;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _tmp_1429 <= _tmp_1428;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _tmp_1430 <= _tmp_1429;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _tmp_1431 <= _tmp_1430;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _tmp_1432 <= _tmp_1431;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _tmp_1433 <= _stream_max_pool_serial_26_source_stop;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _tmp_1434 <= _tmp_1433;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _tmp_1435 <= _tmp_1434;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _tmp_1436 <= _tmp_1435;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _tmp_1437 <= _tmp_1436;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _tmp_1438 <= _tmp_1437;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _tmp_1439 <= _tmp_1438;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _tmp_1440 <= _stream_max_pool_serial_26_source_busy;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _tmp_1441 <= _tmp_1440;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _tmp_1442 <= _tmp_1441;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _tmp_1443 <= _tmp_1442;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _tmp_1444 <= _tmp_1443;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _tmp_1445 <= _tmp_1444;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _tmp_1446 <= _tmp_1445;
      end 
      if(_stream_max_pool_serial_26_stream_oready) begin
        _tmp_1447 <= _stream_max_pool_serial_26_sink_busy;
      end 
      if(!_stream_max_pool_serial_26_sink_busy && _tmp_1447) begin
        _stream_max_pool_serial_26_busy_reg <= 0;
      end 
      if(_stream_max_pool_serial_26_source_busy) begin
        _stream_max_pool_serial_26_busy_reg <= 1;
      end 
    end
  end

  localparam _stream_max_pool_serial_26_fsm_1 = 1;
  localparam _stream_max_pool_serial_26_fsm_2 = 2;
  localparam _stream_max_pool_serial_26_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_max_pool_serial_26_fsm <= _stream_max_pool_serial_26_fsm_init;
      _stream_max_pool_serial_26_source_start <= 0;
      _stream_max_pool_serial_26_source_busy <= 0;
      _stream_max_pool_serial_26_stream_ivalid <= 0;
    end else begin
      if(_stream_max_pool_serial_26_stream_oready && _tmp_1412) begin
        _stream_max_pool_serial_26_stream_ivalid <= 1;
      end 
      if(_stream_max_pool_serial_26_stream_oready && _tmp_1422) begin
        _stream_max_pool_serial_26_stream_ivalid <= 0;
      end 
      case(_stream_max_pool_serial_26_fsm)
        _stream_max_pool_serial_26_fsm_init: begin
          if(_stream_max_pool_serial_26_run_flag) begin
            _stream_max_pool_serial_26_source_start <= 1;
          end 
          if(_stream_max_pool_serial_26_run_flag) begin
            _stream_max_pool_serial_26_fsm <= _stream_max_pool_serial_26_fsm_1;
          end 
        end
        _stream_max_pool_serial_26_fsm_1: begin
          if(_stream_max_pool_serial_26_source_start && _stream_max_pool_serial_26_stream_oready) begin
            _stream_max_pool_serial_26_source_start <= 0;
            _stream_max_pool_serial_26_source_busy <= 1;
          end 
          if(_stream_max_pool_serial_26_source_start && _stream_max_pool_serial_26_stream_oready) begin
            _stream_max_pool_serial_26_fsm <= _stream_max_pool_serial_26_fsm_2;
          end 
        end
        _stream_max_pool_serial_26_fsm_2: begin
          if(_stream_max_pool_serial_26_stream_oready) begin
            _stream_max_pool_serial_26_fsm <= _stream_max_pool_serial_26_fsm_3;
          end 
        end
        _stream_max_pool_serial_26_fsm_3: begin
          if(_stream_max_pool_serial_26_stream_oready && (_stream_max_pool_serial_26_source_1_idle && (_stream_max_pool_serial_26_fsm == 3))) begin
            _stream_max_pool_serial_26_source_busy <= 0;
          end 
          if(_stream_max_pool_serial_26_stream_oready && (_stream_max_pool_serial_26_source_1_idle && (_stream_max_pool_serial_26_fsm == 3)) && _stream_max_pool_serial_26_run_flag) begin
            _stream_max_pool_serial_26_source_start <= 1;
          end 
          if(_stream_max_pool_serial_26_stream_oready && (_stream_max_pool_serial_26_source_1_idle && (_stream_max_pool_serial_26_fsm == 3))) begin
            _stream_max_pool_serial_26_fsm <= _stream_max_pool_serial_26_fsm_init;
          end 
          if(_stream_max_pool_serial_26_stream_oready && (_stream_max_pool_serial_26_source_1_idle && (_stream_max_pool_serial_26_fsm == 3)) && _stream_max_pool_serial_26_run_flag) begin
            _stream_max_pool_serial_26_fsm <= _stream_max_pool_serial_26_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _stream_avg_pool_serial_52_source_1_source_ram_renable <= 0;
      _stream_avg_pool_serial_52_source_1_source_fifo_deq <= 0;
      _stream_avg_pool_serial_52_source_1_idle <= 1;
      _stream_avg_pool_serial_52_sink_5_sink_wenable <= 0;
      _stream_avg_pool_serial_52_sink_5_sink_fifo_enq <= 0;
      _stream_avg_pool_serial_52_sink_6_sink_wenable <= 0;
      _stream_avg_pool_serial_52_sink_6_sink_fifo_enq <= 0;
      __stream_avg_pool_serial_52_stream_ivalid_1 <= 0;
      __stream_avg_pool_serial_52_stream_ivalid_2 <= 0;
      __stream_avg_pool_serial_52_stream_ivalid_3 <= 0;
      __stream_avg_pool_serial_52_stream_ivalid_4 <= 0;
      __stream_avg_pool_serial_52_stream_ivalid_5 <= 0;
      __stream_avg_pool_serial_52_stream_ivalid_6 <= 0;
      _counter_data_916 <= 1'sd0;
      _counter_count_916 <= 1'sd0;
      __delay_data_1183__variable_914 <= 0;
      __delay_data_1184_reinterpretcast_924 <= 0;
      __delay_data_1186__variable_915 <= 0;
      __delay_data_1189__variable_912 <= 0;
      _pointer_data_919 <= 0;
      __delay_data_1185__delay_1184_reinterpretcast_924 <= 0;
      __delay_data_1187__delay_1186__variable_915 <= 0;
      __delay_data_1190__delay_1189__variable_912 <= 0;
      _cond_data_926 <= 0;
      __delay_data_1188__delay_1187__delay_1186__variable_915 <= 0;
      __delay_data_1191__delay_1190__delay_1189__variable_912 <= 0;
      _stream_avg_pool_serial_52_parameter_0_next_parameter_data <= 0;
      __variable_wdata_912 <= 0;
      _stream_avg_pool_serial_52_parameter_2_next_parameter_data <= 0;
      __variable_wdata_914 <= 0;
      _stream_avg_pool_serial_52_source_1_source_mode <= 5'b0;
      _stream_avg_pool_serial_52_source_1_source_offset <= 0;
      _source_stream_avg_pool_serial_52_source_1_pat_size_0 <= 0;
      _source_stream_avg_pool_serial_52_source_1_pat_stride_0 <= 0;
      _source_stream_avg_pool_serial_52_source_1_pat_size_1 <= 0;
      _source_stream_avg_pool_serial_52_source_1_pat_stride_1 <= 0;
      _source_stream_avg_pool_serial_52_source_1_pat_size_2 <= 0;
      _source_stream_avg_pool_serial_52_source_1_pat_stride_2 <= 0;
      _source_stream_avg_pool_serial_52_source_1_pat_size_3 <= 0;
      _source_stream_avg_pool_serial_52_source_1_pat_stride_3 <= 0;
      _stream_avg_pool_serial_52_source_1_source_sel <= 0;
      _stream_avg_pool_serial_52_source_1_source_offset_buf <= 0;
      _source_stream_avg_pool_serial_52_source_1_pat_cur_offset_0 <= 0;
      _source_stream_avg_pool_serial_52_source_1_pat_cur_offset_1 <= 0;
      _source_stream_avg_pool_serial_52_source_1_pat_cur_offset_2 <= 0;
      _source_stream_avg_pool_serial_52_source_1_pat_cur_offset_3 <= 0;
      _source_stream_avg_pool_serial_52_source_1_pat_count_0 <= 0;
      _source_stream_avg_pool_serial_52_source_1_pat_count_1 <= 0;
      _source_stream_avg_pool_serial_52_source_1_pat_count_2 <= 0;
      _source_stream_avg_pool_serial_52_source_1_pat_count_3 <= 0;
      _source_stream_avg_pool_serial_52_source_1_pat_size_buf_0 <= 0;
      _source_stream_avg_pool_serial_52_source_1_pat_size_buf_1 <= 0;
      _source_stream_avg_pool_serial_52_source_1_pat_size_buf_2 <= 0;
      _source_stream_avg_pool_serial_52_source_1_pat_size_buf_3 <= 0;
      _source_stream_avg_pool_serial_52_source_1_pat_stride_buf_0 <= 0;
      _source_stream_avg_pool_serial_52_source_1_pat_stride_buf_1 <= 0;
      _source_stream_avg_pool_serial_52_source_1_pat_stride_buf_2 <= 0;
      _source_stream_avg_pool_serial_52_source_1_pat_stride_buf_3 <= 0;
      __variable_wdata_913 <= 0;
      _stream_avg_pool_serial_52_source_1_source_ram_raddr <= 0;
      _tmp_1508 <= 0;
      _tmp_1509 <= 0;
      _tmp_1510 <= 0;
      _tmp_1511 <= 0;
      _tmp_1512 <= 0;
      _tmp_1513 <= 0;
      _tmp_1514 <= 0;
      _tmp_1515 <= 0;
      _tmp_1518 <= 0;
      _tmp_1519 <= 0;
      _tmp_1520 <= 0;
      _tmp_1521 <= 0;
      _tmp_1522 <= 0;
      _tmp_1523 <= 0;
      _tmp_1524 <= 0;
      _tmp_1525 <= 0;
      _tmp_1526 <= 0;
      _tmp_1527 <= 0;
      _tmp_1528 <= 0;
      _tmp_1529 <= 0;
      _tmp_1530 <= 0;
      _tmp_1531 <= 0;
      _tmp_1532 <= 0;
      _tmp_1533 <= 0;
      _stream_avg_pool_serial_52_sink_5_sink_mode <= 5'b0;
      _stream_avg_pool_serial_52_sink_5_sink_offset <= 0;
      _stream_avg_pool_serial_52_sink_5_sink_size <= 0;
      _stream_avg_pool_serial_52_sink_5_sink_stride <= 0;
      _stream_avg_pool_serial_52_sink_5_sink_sel <= 0;
      _stream_avg_pool_serial_52_sink_5_sink_offset_buf <= 0;
      _stream_avg_pool_serial_52_sink_5_sink_size_buf <= 0;
      _stream_avg_pool_serial_52_sink_5_sink_stride_buf <= 0;
      _stream_avg_pool_serial_52_sink_5_sink_waddr <= 0;
      _stream_avg_pool_serial_52_sink_5_sink_count <= 0;
      _stream_avg_pool_serial_52_sink_5_sink_wdata <= 0;
      _tmp_1559 <= 0;
      _tmp_1560 <= 0;
      _tmp_1561 <= 0;
      _tmp_1562 <= 0;
      _tmp_1563 <= 0;
      _tmp_1564 <= 0;
      __variable_wdata_915 <= 0;
      _tmp_1565 <= 0;
      _tmp_1566 <= 0;
      _tmp_1567 <= 0;
      _tmp_1568 <= 0;
      _tmp_1571 <= 0;
      _tmp_1574 <= 0;
      _tmp_1575 <= 0;
      _tmp_1576 <= 0;
      _tmp_1577 <= 0;
      _tmp_1578 <= 0;
      _tmp_1579 <= 0;
      _tmp_1580 <= 0;
      _tmp_1581 <= 0;
      _tmp_1582 <= 0;
      _tmp_1583 <= 0;
      _tmp_1584 <= 0;
      _tmp_1585 <= 0;
      _tmp_1586 <= 0;
      _tmp_1587 <= 0;
      _tmp_1588 <= 0;
      _tmp_1589 <= 0;
      _tmp_1590 <= 0;
      _tmp_1591 <= 0;
      _tmp_1592 <= 0;
      _tmp_1593 <= 0;
      _tmp_1594 <= 0;
      _tmp_1595 <= 0;
      _tmp_1596 <= 0;
      _tmp_1597 <= 0;
      _tmp_1598 <= 0;
      _tmp_1599 <= 0;
      _stream_avg_pool_serial_52_busy_reg <= 0;
    end else begin
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _stream_avg_pool_serial_52_source_1_source_ram_renable <= 0;
        _stream_avg_pool_serial_52_source_1_source_fifo_deq <= 0;
      end 
      _stream_avg_pool_serial_52_source_1_idle <= _stream_avg_pool_serial_52_source_1_idle;
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _stream_avg_pool_serial_52_sink_5_sink_wenable <= 0;
        _stream_avg_pool_serial_52_sink_5_sink_fifo_enq <= 0;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _stream_avg_pool_serial_52_sink_6_sink_wenable <= 0;
        _stream_avg_pool_serial_52_sink_6_sink_fifo_enq <= 0;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        __stream_avg_pool_serial_52_stream_ivalid_1 <= _stream_avg_pool_serial_52_stream_ivalid;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        __stream_avg_pool_serial_52_stream_ivalid_2 <= __stream_avg_pool_serial_52_stream_ivalid_1;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        __stream_avg_pool_serial_52_stream_ivalid_3 <= __stream_avg_pool_serial_52_stream_ivalid_2;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        __stream_avg_pool_serial_52_stream_ivalid_4 <= __stream_avg_pool_serial_52_stream_ivalid_3;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        __stream_avg_pool_serial_52_stream_ivalid_5 <= __stream_avg_pool_serial_52_stream_ivalid_4;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        __stream_avg_pool_serial_52_stream_ivalid_6 <= __stream_avg_pool_serial_52_stream_ivalid_5;
      end 
      if(_stream_avg_pool_serial_52_stream_ivalid && _stream_avg_pool_serial_52_stream_oready && _counter_reset_cond_916) begin
        _counter_data_916 <= 1'sd0;
      end 
      if(_stream_avg_pool_serial_52_stream_ivalid && _stream_avg_pool_serial_52_stream_oready) begin
        _counter_data_916 <= _counter_current_count_916;
      end 
      if(_stream_avg_pool_serial_52_stream_ivalid && _stream_avg_pool_serial_52_stream_oready) begin
        _counter_count_916 <= (_counter_current_count_916 >= stream_avg_pool_serial_52_parameter_0_data - 2'sd1)? _counter_current_count_916 + 2'sd1 - stream_avg_pool_serial_52_parameter_0_data : _counter_current_count_916 + 2'sd1;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        __delay_data_1183__variable_914 <= stream_avg_pool_serial_52_parameter_2_data;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        __delay_data_1184_reinterpretcast_924 <= _reinterpretcast_data_924;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        __delay_data_1186__variable_915 <= stream_avg_pool_serial_52__reduce_reset_data;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        __delay_data_1189__variable_912 <= stream_avg_pool_serial_52_parameter_0_data;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _pointer_data_919 <= __delay_data_1183__variable_914[_counter_data_916];
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        __delay_data_1185__delay_1184_reinterpretcast_924 <= __delay_data_1184_reinterpretcast_924;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        __delay_data_1187__delay_1186__variable_915 <= __delay_data_1186__variable_915;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        __delay_data_1190__delay_1189__variable_912 <= __delay_data_1189__variable_912;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _cond_data_926 <= (_pointer_data_919)? 1'sd0 : __delay_data_1185__delay_1184_reinterpretcast_924;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        __delay_data_1188__delay_1187__delay_1186__variable_915 <= __delay_data_1187__delay_1186__variable_915;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        __delay_data_1191__delay_1190__delay_1189__variable_912 <= __delay_data_1190__delay_1189__variable_912;
      end 
      if(_set_flag_1492) begin
        _stream_avg_pool_serial_52_parameter_0_next_parameter_data <= 1;
      end 
      if(_stream_avg_pool_serial_52_source_start) begin
        __variable_wdata_912 <= _stream_avg_pool_serial_52_parameter_0_next_parameter_data;
      end 
      if(_set_flag_1493) begin
        _stream_avg_pool_serial_52_parameter_2_next_parameter_data <= avg_pool_serial_52_stream_pad_masks;
      end 
      if(_stream_avg_pool_serial_52_source_start) begin
        __variable_wdata_914 <= _stream_avg_pool_serial_52_parameter_2_next_parameter_data;
      end 
      if(_set_flag_1494) begin
        _stream_avg_pool_serial_52_source_1_source_mode <= 5'b10;
        _stream_avg_pool_serial_52_source_1_source_offset <= avg_pool_serial_52_stream_act_local + avg_pool_serial_52_act_page_comp_offset_buf;
      end 
      if(_set_flag_1494) begin
        _source_stream_avg_pool_serial_52_source_1_pat_size_0 <= 1;
        _source_stream_avg_pool_serial_52_source_1_pat_stride_0 <= cparam_avg_pool_serial_52_act_read_block;
      end 
      if(_set_flag_1494) begin
        _source_stream_avg_pool_serial_52_source_1_pat_size_1 <= 1;
        _source_stream_avg_pool_serial_52_source_1_pat_stride_1 <= cparam_avg_pool_serial_52_act_read_size;
      end 
      if(_set_flag_1494) begin
        _source_stream_avg_pool_serial_52_source_1_pat_size_2 <= cparam_avg_pool_serial_52_stream_size;
        _source_stream_avg_pool_serial_52_source_1_pat_stride_2 <= 1;
      end 
      if(_set_flag_1494) begin
        _source_stream_avg_pool_serial_52_source_1_pat_size_3 <= 1;
        _source_stream_avg_pool_serial_52_source_1_pat_stride_3 <= 0;
      end 
      if(_set_flag_1494) begin
        _stream_avg_pool_serial_52_source_1_source_sel <= 1;
      end 
      if(_stream_avg_pool_serial_52_source_start && _stream_avg_pool_serial_52_source_1_source_mode & 5'b10 && _stream_avg_pool_serial_52_stream_oready) begin
        _stream_avg_pool_serial_52_source_1_source_offset_buf <= _stream_avg_pool_serial_52_source_1_source_offset;
      end 
      if(_stream_avg_pool_serial_52_source_start && _stream_avg_pool_serial_52_source_1_source_mode & 5'b10 && _stream_avg_pool_serial_52_stream_oready) begin
        _source_stream_avg_pool_serial_52_source_1_pat_cur_offset_0 <= 0;
      end 
      if(_stream_avg_pool_serial_52_source_start && _stream_avg_pool_serial_52_source_1_source_mode & 5'b10 && _stream_avg_pool_serial_52_stream_oready) begin
        _source_stream_avg_pool_serial_52_source_1_pat_cur_offset_1 <= 0;
      end 
      if(_stream_avg_pool_serial_52_source_start && _stream_avg_pool_serial_52_source_1_source_mode & 5'b10 && _stream_avg_pool_serial_52_stream_oready) begin
        _source_stream_avg_pool_serial_52_source_1_pat_cur_offset_2 <= 0;
      end 
      if(_stream_avg_pool_serial_52_source_start && _stream_avg_pool_serial_52_source_1_source_mode & 5'b10 && _stream_avg_pool_serial_52_stream_oready) begin
        _source_stream_avg_pool_serial_52_source_1_pat_cur_offset_3 <= 0;
      end 
      if(_stream_avg_pool_serial_52_source_start && _stream_avg_pool_serial_52_source_1_source_mode & 5'b10 && _stream_avg_pool_serial_52_stream_oready) begin
        _source_stream_avg_pool_serial_52_source_1_pat_count_0 <= _source_stream_avg_pool_serial_52_source_1_pat_size_0 - 1;
      end 
      if(_stream_avg_pool_serial_52_source_start && _stream_avg_pool_serial_52_source_1_source_mode & 5'b10 && _stream_avg_pool_serial_52_stream_oready) begin
        _source_stream_avg_pool_serial_52_source_1_pat_count_1 <= _source_stream_avg_pool_serial_52_source_1_pat_size_1 - 1;
      end 
      if(_stream_avg_pool_serial_52_source_start && _stream_avg_pool_serial_52_source_1_source_mode & 5'b10 && _stream_avg_pool_serial_52_stream_oready) begin
        _source_stream_avg_pool_serial_52_source_1_pat_count_2 <= _source_stream_avg_pool_serial_52_source_1_pat_size_2 - 1;
      end 
      if(_stream_avg_pool_serial_52_source_start && _stream_avg_pool_serial_52_source_1_source_mode & 5'b10 && _stream_avg_pool_serial_52_stream_oready) begin
        _source_stream_avg_pool_serial_52_source_1_pat_count_3 <= _source_stream_avg_pool_serial_52_source_1_pat_size_3 - 1;
      end 
      if(_stream_avg_pool_serial_52_source_start && _stream_avg_pool_serial_52_source_1_source_mode & 5'b10 && _stream_avg_pool_serial_52_stream_oready) begin
        _source_stream_avg_pool_serial_52_source_1_pat_size_buf_0 <= _source_stream_avg_pool_serial_52_source_1_pat_size_0;
      end 
      if(_stream_avg_pool_serial_52_source_start && _stream_avg_pool_serial_52_source_1_source_mode & 5'b10 && _stream_avg_pool_serial_52_stream_oready) begin
        _source_stream_avg_pool_serial_52_source_1_pat_size_buf_1 <= _source_stream_avg_pool_serial_52_source_1_pat_size_1;
      end 
      if(_stream_avg_pool_serial_52_source_start && _stream_avg_pool_serial_52_source_1_source_mode & 5'b10 && _stream_avg_pool_serial_52_stream_oready) begin
        _source_stream_avg_pool_serial_52_source_1_pat_size_buf_2 <= _source_stream_avg_pool_serial_52_source_1_pat_size_2;
      end 
      if(_stream_avg_pool_serial_52_source_start && _stream_avg_pool_serial_52_source_1_source_mode & 5'b10 && _stream_avg_pool_serial_52_stream_oready) begin
        _source_stream_avg_pool_serial_52_source_1_pat_size_buf_3 <= _source_stream_avg_pool_serial_52_source_1_pat_size_3;
      end 
      if(_stream_avg_pool_serial_52_source_start && _stream_avg_pool_serial_52_source_1_source_mode & 5'b10 && _stream_avg_pool_serial_52_stream_oready) begin
        _source_stream_avg_pool_serial_52_source_1_pat_stride_buf_0 <= _source_stream_avg_pool_serial_52_source_1_pat_stride_0;
      end 
      if(_stream_avg_pool_serial_52_source_start && _stream_avg_pool_serial_52_source_1_source_mode & 5'b10 && _stream_avg_pool_serial_52_stream_oready) begin
        _source_stream_avg_pool_serial_52_source_1_pat_stride_buf_1 <= _source_stream_avg_pool_serial_52_source_1_pat_stride_1;
      end 
      if(_stream_avg_pool_serial_52_source_start && _stream_avg_pool_serial_52_source_1_source_mode & 5'b10 && _stream_avg_pool_serial_52_stream_oready) begin
        _source_stream_avg_pool_serial_52_source_1_pat_stride_buf_2 <= _source_stream_avg_pool_serial_52_source_1_pat_stride_2;
      end 
      if(_stream_avg_pool_serial_52_source_start && _stream_avg_pool_serial_52_source_1_source_mode & 5'b10 && _stream_avg_pool_serial_52_stream_oready) begin
        _source_stream_avg_pool_serial_52_source_1_pat_stride_buf_3 <= _source_stream_avg_pool_serial_52_source_1_pat_stride_3;
      end 
      if(_stream_avg_pool_serial_52_stream_oready && _stream_avg_pool_serial_52_source_busy && _stream_avg_pool_serial_52_is_root) begin
        __variable_wdata_913 <= _stream_avg_pool_serial_52_source_1_source_ram_rdata;
      end 
      if((_stream_avg_pool_serial_52_source_1_source_pat_fsm_0 == 1) && _stream_avg_pool_serial_52_stream_oready) begin
        _stream_avg_pool_serial_52_source_1_idle <= 0;
        _stream_avg_pool_serial_52_source_1_source_ram_raddr <= _stream_avg_pool_serial_52_source_1_source_pat_all_offset;
        _stream_avg_pool_serial_52_source_1_source_ram_renable <= 1;
      end 
      if((_stream_avg_pool_serial_52_source_1_source_pat_fsm_0 == 1) && _stream_avg_pool_serial_52_stream_oready) begin
        _source_stream_avg_pool_serial_52_source_1_pat_cur_offset_0 <= _source_stream_avg_pool_serial_52_source_1_pat_cur_offset_0 + _source_stream_avg_pool_serial_52_source_1_pat_stride_buf_0;
        _source_stream_avg_pool_serial_52_source_1_pat_count_0 <= _source_stream_avg_pool_serial_52_source_1_pat_count_0 - 1;
      end 
      if((_stream_avg_pool_serial_52_source_1_source_pat_fsm_0 == 1) && (_source_stream_avg_pool_serial_52_source_1_pat_count_0 == 0) && _stream_avg_pool_serial_52_stream_oready) begin
        _source_stream_avg_pool_serial_52_source_1_pat_cur_offset_0 <= 0;
        _source_stream_avg_pool_serial_52_source_1_pat_count_0 <= _source_stream_avg_pool_serial_52_source_1_pat_size_buf_0 - 1;
      end 
      if((_stream_avg_pool_serial_52_source_1_source_pat_fsm_0 == 1) && (_source_stream_avg_pool_serial_52_source_1_pat_count_0 == 0) && _stream_avg_pool_serial_52_stream_oready) begin
        _source_stream_avg_pool_serial_52_source_1_pat_cur_offset_1 <= _source_stream_avg_pool_serial_52_source_1_pat_cur_offset_1 + _source_stream_avg_pool_serial_52_source_1_pat_stride_buf_1;
        _source_stream_avg_pool_serial_52_source_1_pat_count_1 <= _source_stream_avg_pool_serial_52_source_1_pat_count_1 - 1;
      end 
      if((_stream_avg_pool_serial_52_source_1_source_pat_fsm_0 == 1) && (_source_stream_avg_pool_serial_52_source_1_pat_count_0 == 0) && (_source_stream_avg_pool_serial_52_source_1_pat_count_1 == 0) && _stream_avg_pool_serial_52_stream_oready) begin
        _source_stream_avg_pool_serial_52_source_1_pat_cur_offset_1 <= 0;
        _source_stream_avg_pool_serial_52_source_1_pat_count_1 <= _source_stream_avg_pool_serial_52_source_1_pat_size_buf_1 - 1;
      end 
      if((_stream_avg_pool_serial_52_source_1_source_pat_fsm_0 == 1) && ((_source_stream_avg_pool_serial_52_source_1_pat_count_0 == 0) && (_source_stream_avg_pool_serial_52_source_1_pat_count_1 == 0)) && _stream_avg_pool_serial_52_stream_oready) begin
        _source_stream_avg_pool_serial_52_source_1_pat_cur_offset_2 <= _source_stream_avg_pool_serial_52_source_1_pat_cur_offset_2 + _source_stream_avg_pool_serial_52_source_1_pat_stride_buf_2;
        _source_stream_avg_pool_serial_52_source_1_pat_count_2 <= _source_stream_avg_pool_serial_52_source_1_pat_count_2 - 1;
      end 
      if((_stream_avg_pool_serial_52_source_1_source_pat_fsm_0 == 1) && ((_source_stream_avg_pool_serial_52_source_1_pat_count_0 == 0) && (_source_stream_avg_pool_serial_52_source_1_pat_count_1 == 0)) && (_source_stream_avg_pool_serial_52_source_1_pat_count_2 == 0) && _stream_avg_pool_serial_52_stream_oready) begin
        _source_stream_avg_pool_serial_52_source_1_pat_cur_offset_2 <= 0;
        _source_stream_avg_pool_serial_52_source_1_pat_count_2 <= _source_stream_avg_pool_serial_52_source_1_pat_size_buf_2 - 1;
      end 
      if((_stream_avg_pool_serial_52_source_1_source_pat_fsm_0 == 1) && ((_source_stream_avg_pool_serial_52_source_1_pat_count_0 == 0) && (_source_stream_avg_pool_serial_52_source_1_pat_count_1 == 0) && (_source_stream_avg_pool_serial_52_source_1_pat_count_2 == 0)) && _stream_avg_pool_serial_52_stream_oready) begin
        _source_stream_avg_pool_serial_52_source_1_pat_cur_offset_3 <= _source_stream_avg_pool_serial_52_source_1_pat_cur_offset_3 + _source_stream_avg_pool_serial_52_source_1_pat_stride_buf_3;
        _source_stream_avg_pool_serial_52_source_1_pat_count_3 <= _source_stream_avg_pool_serial_52_source_1_pat_count_3 - 1;
      end 
      if((_stream_avg_pool_serial_52_source_1_source_pat_fsm_0 == 1) && ((_source_stream_avg_pool_serial_52_source_1_pat_count_0 == 0) && (_source_stream_avg_pool_serial_52_source_1_pat_count_1 == 0) && (_source_stream_avg_pool_serial_52_source_1_pat_count_2 == 0)) && (_source_stream_avg_pool_serial_52_source_1_pat_count_3 == 0) && _stream_avg_pool_serial_52_stream_oready) begin
        _source_stream_avg_pool_serial_52_source_1_pat_cur_offset_3 <= 0;
        _source_stream_avg_pool_serial_52_source_1_pat_count_3 <= _source_stream_avg_pool_serial_52_source_1_pat_size_buf_3 - 1;
      end 
      if((_stream_avg_pool_serial_52_source_1_source_pat_fsm_0 == 1) && _stream_avg_pool_serial_52_source_stop && _stream_avg_pool_serial_52_stream_oready) begin
        _stream_avg_pool_serial_52_source_1_source_ram_renable <= 0;
        _stream_avg_pool_serial_52_source_1_idle <= 1;
      end 
      if((_stream_avg_pool_serial_52_source_1_source_pat_fsm_0 == 2) && _stream_avg_pool_serial_52_stream_oready) begin
        _stream_avg_pool_serial_52_source_1_source_ram_renable <= 0;
        _stream_avg_pool_serial_52_source_1_idle <= 1;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1508 <= _set_flag_1507;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1509 <= _tmp_1508;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1510 <= _tmp_1509;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1511 <= _tmp_1510;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1512 <= _tmp_1511;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1513 <= _tmp_1512;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1514 <= _tmp_1513;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1515 <= _tmp_1514;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1518 <= _tmp_1517;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1519 <= _tmp_1518;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1520 <= _tmp_1519;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1521 <= _tmp_1520;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1522 <= _tmp_1521;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1523 <= _tmp_1522;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1524 <= _tmp_1523;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1525 <= _tmp_1524;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1526 <= cparam_avg_pool_serial_52_stream_size;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1527 <= _tmp_1526;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1528 <= _tmp_1527;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1529 <= _tmp_1528;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1530 <= _tmp_1529;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1531 <= _tmp_1530;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1532 <= _tmp_1531;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1533 <= _tmp_1532;
      end 
      if(_tmp_1515) begin
        _stream_avg_pool_serial_52_sink_5_sink_mode <= 5'b1;
        _stream_avg_pool_serial_52_sink_5_sink_offset <= _tmp_1525;
        _stream_avg_pool_serial_52_sink_5_sink_size <= _tmp_1533;
        _stream_avg_pool_serial_52_sink_5_sink_stride <= 1;
      end 
      if(_tmp_1515) begin
        _stream_avg_pool_serial_52_sink_5_sink_sel <= 2;
      end 
      if(_stream_avg_pool_serial_52_sink_start && _stream_avg_pool_serial_52_sink_5_sink_mode & 5'b1 && _stream_avg_pool_serial_52_stream_oready) begin
        _stream_avg_pool_serial_52_sink_5_sink_offset_buf <= _stream_avg_pool_serial_52_sink_5_sink_offset;
        _stream_avg_pool_serial_52_sink_5_sink_size_buf <= _stream_avg_pool_serial_52_sink_5_sink_size;
        _stream_avg_pool_serial_52_sink_5_sink_stride_buf <= _stream_avg_pool_serial_52_sink_5_sink_stride;
      end 
      if((_stream_avg_pool_serial_52_sink_5_sink_fsm_1 == 1) && _stream_avg_pool_serial_52_stream_oready) begin
        _stream_avg_pool_serial_52_sink_5_sink_waddr <= _stream_avg_pool_serial_52_sink_5_sink_offset_buf - _stream_avg_pool_serial_52_sink_5_sink_stride_buf;
        _stream_avg_pool_serial_52_sink_5_sink_count <= _stream_avg_pool_serial_52_sink_5_sink_size_buf;
      end 
      if((_stream_avg_pool_serial_52_sink_5_sink_fsm_1 == 2) && stream_avg_pool_serial_52_sink_6_data && _stream_avg_pool_serial_52_stream_oready) begin
        _stream_avg_pool_serial_52_sink_5_sink_waddr <= _stream_avg_pool_serial_52_sink_5_sink_waddr + _stream_avg_pool_serial_52_sink_5_sink_stride_buf;
        _stream_avg_pool_serial_52_sink_5_sink_wdata <= stream_avg_pool_serial_52_sink_5_data;
        _stream_avg_pool_serial_52_sink_5_sink_wenable <= 1;
        _stream_avg_pool_serial_52_sink_5_sink_count <= _stream_avg_pool_serial_52_sink_5_sink_count - 1;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1559 <= _stream_avg_pool_serial_52_source_start;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1560 <= _tmp_1559;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1561 <= _tmp_1560;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1562 <= _stream_avg_pool_serial_52_source_start;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1563 <= _tmp_1562;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1564 <= _tmp_1563;
      end 
      if(_stream_avg_pool_serial_52_stream_oready && _tmp_1564) begin
        __variable_wdata_915 <= 1;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1565 <= _stream_avg_pool_serial_52_source_start;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1566 <= _tmp_1565;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1567 <= _tmp_1566;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1568 <= _tmp_1567;
      end 
      if(_stream_avg_pool_serial_52_stream_oready && _tmp_1568) begin
        __variable_wdata_915 <= 0;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1571 <= _tmp_1570;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1574 <= _tmp_1573;
      end 
      if(_stream_avg_pool_serial_52_stream_oready && _tmp_1574) begin
        __variable_wdata_915 <= 1;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1575 <= _stream_avg_pool_serial_52_source_start;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1576 <= _tmp_1575;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1577 <= _tmp_1576;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1578 <= _tmp_1577;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1579 <= _tmp_1578;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1580 <= _tmp_1579;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1581 <= _tmp_1580;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1582 <= _tmp_1581;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1583 <= _stream_avg_pool_serial_52_source_stop;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1584 <= _tmp_1583;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1585 <= _tmp_1584;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1586 <= _tmp_1585;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1587 <= _tmp_1586;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1588 <= _tmp_1587;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1589 <= _tmp_1588;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1590 <= _tmp_1589;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1591 <= _stream_avg_pool_serial_52_source_busy;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1592 <= _tmp_1591;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1593 <= _tmp_1592;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1594 <= _tmp_1593;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1595 <= _tmp_1594;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1596 <= _tmp_1595;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1597 <= _tmp_1596;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1598 <= _tmp_1597;
      end 
      if(_stream_avg_pool_serial_52_stream_oready) begin
        _tmp_1599 <= _stream_avg_pool_serial_52_sink_busy;
      end 
      if(!_stream_avg_pool_serial_52_sink_busy && _tmp_1599) begin
        _stream_avg_pool_serial_52_busy_reg <= 0;
      end 
      if(_stream_avg_pool_serial_52_source_busy) begin
        _stream_avg_pool_serial_52_busy_reg <= 1;
      end 
    end
  end

  localparam _stream_avg_pool_serial_52_fsm_1 = 1;
  localparam _stream_avg_pool_serial_52_fsm_2 = 2;
  localparam _stream_avg_pool_serial_52_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_avg_pool_serial_52_fsm <= _stream_avg_pool_serial_52_fsm_init;
      _stream_avg_pool_serial_52_source_start <= 0;
      _stream_avg_pool_serial_52_source_busy <= 0;
      _stream_avg_pool_serial_52_stream_ivalid <= 0;
    end else begin
      if(_stream_avg_pool_serial_52_stream_oready && _tmp_1561) begin
        _stream_avg_pool_serial_52_stream_ivalid <= 1;
      end 
      if(_stream_avg_pool_serial_52_stream_oready && _tmp_1571) begin
        _stream_avg_pool_serial_52_stream_ivalid <= 0;
      end 
      case(_stream_avg_pool_serial_52_fsm)
        _stream_avg_pool_serial_52_fsm_init: begin
          if(_stream_avg_pool_serial_52_run_flag) begin
            _stream_avg_pool_serial_52_source_start <= 1;
          end 
          if(_stream_avg_pool_serial_52_run_flag) begin
            _stream_avg_pool_serial_52_fsm <= _stream_avg_pool_serial_52_fsm_1;
          end 
        end
        _stream_avg_pool_serial_52_fsm_1: begin
          if(_stream_avg_pool_serial_52_source_start && _stream_avg_pool_serial_52_stream_oready) begin
            _stream_avg_pool_serial_52_source_start <= 0;
            _stream_avg_pool_serial_52_source_busy <= 1;
          end 
          if(_stream_avg_pool_serial_52_source_start && _stream_avg_pool_serial_52_stream_oready) begin
            _stream_avg_pool_serial_52_fsm <= _stream_avg_pool_serial_52_fsm_2;
          end 
        end
        _stream_avg_pool_serial_52_fsm_2: begin
          if(_stream_avg_pool_serial_52_stream_oready) begin
            _stream_avg_pool_serial_52_fsm <= _stream_avg_pool_serial_52_fsm_3;
          end 
        end
        _stream_avg_pool_serial_52_fsm_3: begin
          if(_stream_avg_pool_serial_52_stream_oready && (_stream_avg_pool_serial_52_source_1_idle && (_stream_avg_pool_serial_52_fsm == 3))) begin
            _stream_avg_pool_serial_52_source_busy <= 0;
          end 
          if(_stream_avg_pool_serial_52_stream_oready && (_stream_avg_pool_serial_52_source_1_idle && (_stream_avg_pool_serial_52_fsm == 3)) && _stream_avg_pool_serial_52_run_flag) begin
            _stream_avg_pool_serial_52_source_start <= 1;
          end 
          if(_stream_avg_pool_serial_52_stream_oready && (_stream_avg_pool_serial_52_source_1_idle && (_stream_avg_pool_serial_52_fsm == 3))) begin
            _stream_avg_pool_serial_52_fsm <= _stream_avg_pool_serial_52_fsm_init;
          end 
          if(_stream_avg_pool_serial_52_stream_oready && (_stream_avg_pool_serial_52_source_1_idle && (_stream_avg_pool_serial_52_fsm == 3)) && _stream_avg_pool_serial_52_run_flag) begin
            _stream_avg_pool_serial_52_fsm <= _stream_avg_pool_serial_52_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _stream_matmul_55_source_7_source_ram_renable <= 0;
      _stream_matmul_55_source_7_source_fifo_deq <= 0;
      _stream_matmul_55_source_7_idle <= 1;
      _stream_matmul_55_source_9_source_ram_renable <= 0;
      _stream_matmul_55_source_9_source_fifo_deq <= 0;
      _stream_matmul_55_source_9_idle <= 1;
      _stream_matmul_55_source_11_source_ram_renable <= 0;
      _stream_matmul_55_source_11_source_fifo_deq <= 0;
      _stream_matmul_55_source_11_idle <= 1;
      _stream_matmul_55_source_13_source_ram_renable <= 0;
      _stream_matmul_55_source_13_source_fifo_deq <= 0;
      _stream_matmul_55_source_13_idle <= 1;
      _stream_matmul_55_source_15_source_ram_renable <= 0;
      _stream_matmul_55_source_15_source_fifo_deq <= 0;
      _stream_matmul_55_source_15_idle <= 1;
      _stream_matmul_55_source_20_source_ram_renable <= 0;
      _stream_matmul_55_source_20_source_fifo_deq <= 0;
      _stream_matmul_55_source_20_idle <= 1;
      _stream_matmul_55_source_21_source_ram_renable <= 0;
      _stream_matmul_55_source_21_source_fifo_deq <= 0;
      _stream_matmul_55_source_21_idle <= 1;
      _stream_matmul_55_sink_26_sink_wenable <= 0;
      _stream_matmul_55_sink_26_sink_fifo_enq <= 0;
      _stream_matmul_55_sink_27_sink_wenable <= 0;
      _stream_matmul_55_sink_27_sink_fifo_enq <= 0;
      __stream_matmul_55_stream_ivalid_1 <= 0;
      __stream_matmul_55_stream_ivalid_2 <= 0;
      __stream_matmul_55_stream_ivalid_3 <= 0;
      __stream_matmul_55_stream_ivalid_4 <= 0;
      __stream_matmul_55_stream_ivalid_5 <= 0;
      __stream_matmul_55_stream_ivalid_6 <= 0;
      __stream_matmul_55_stream_ivalid_7 <= 0;
      __stream_matmul_55_stream_ivalid_8 <= 0;
      __stream_matmul_55_stream_ivalid_9 <= 0;
      __stream_matmul_55_stream_ivalid_10 <= 0;
      __stream_matmul_55_stream_ivalid_11 <= 0;
      __stream_matmul_55_stream_ivalid_12 <= 0;
      __stream_matmul_55_stream_ivalid_13 <= 0;
      __stream_matmul_55_stream_ivalid_14 <= 0;
      __stream_matmul_55_stream_ivalid_15 <= 0;
      __stream_matmul_55_stream_ivalid_16 <= 0;
      __stream_matmul_55_stream_ivalid_17 <= 0;
      __stream_matmul_55_stream_ivalid_18 <= 0;
      __stream_matmul_55_stream_ivalid_19 <= 0;
      __stream_matmul_55_stream_ivalid_20 <= 0;
      __stream_matmul_55_stream_ivalid_21 <= 0;
      __stream_matmul_55_stream_ivalid_22 <= 0;
      __stream_matmul_55_stream_ivalid_23 <= 0;
      __stream_matmul_55_stream_ivalid_24 <= 0;
      __stream_matmul_55_stream_ivalid_25 <= 0;
      __stream_matmul_55_stream_ivalid_26 <= 0;
      __stream_matmul_55_stream_ivalid_27 <= 0;
      __stream_matmul_55_stream_ivalid_28 <= 0;
      __stream_matmul_55_stream_ivalid_29 <= 0;
      _eq_data_991 <= 0;
      _eq_data_995 <= 0;
      _plus_data_1015 <= 0;
      _plus_data_1020 <= 0;
      _plus_data_1025 <= 0;
      _eq_data_1031 <= 0;
      _eq_data_1034 <= 0;
      __delay_data_1192__variable_990 <= 0;
      __delay_data_1193_pointer_1010 <= 0;
      __delay_data_1194_reinterpretcast_1009 <= 0;
      __delay_data_1195__variable_941 <= 0;
      __delay_data_1216__variable_936 <= 0;
      __delay_data_1227_cond_957 <= 0;
      __delay_data_1244_cond_964 <= 0;
      __delay_data_1196__delay_1195__variable_941 <= 0;
      __delay_data_1206_plus_1020 <= 0;
      __delay_data_1217__delay_1216__variable_936 <= 0;
      __delay_data_1228__delay_1227_cond_957 <= 0;
      __delay_data_1245__delay_1244_cond_964 <= 0;
      __delay_data_1262_plus_1025 <= 0;
      __delay_data_1280_eq_1031 <= 0;
      __delay_data_1309_eq_1034 <= 0;
      __delay_data_1197__delay_1196__delay_1195__variable_941 <= 0;
      __delay_data_1207__delay_1206_plus_1020 <= 0;
      __delay_data_1218__delay_1217__delay_1216__variable_936 <= 0;
      __delay_data_1229__delay_1228__delay_1227_cond_957 <= 0;
      __delay_data_1246__delay_1245__delay_1244_cond_964 <= 0;
      __delay_data_1263__delay_1262_plus_1025 <= 0;
      __delay_data_1281__delay_1280_eq_1031 <= 0;
      __delay_data_1310__delay_1309_eq_1034 <= 0;
      __delay_data_1198__delay_1197__delay_1196____variable_941 <= 0;
      __delay_data_1208__delay_1207__delay_1206_plus_1020 <= 0;
      __delay_data_1219__delay_1218__delay_1217____variable_936 <= 0;
      __delay_data_1230__delay_1229__delay_1228__delay_1227_cond_957 <= 0;
      __delay_data_1247__delay_1246__delay_1245__delay_1244_cond_964 <= 0;
      __delay_data_1264__delay_1263__delay_1262_plus_1025 <= 0;
      __delay_data_1282__delay_1281__delay_1280_eq_1031 <= 0;
      __delay_data_1311__delay_1310__delay_1309_eq_1034 <= 0;
      __delay_data_1199__delay_1198__delay_1197____variable_941 <= 0;
      __delay_data_1209__delay_1208__delay_1207___plus_1020 <= 0;
      __delay_data_1220__delay_1219__delay_1218____variable_936 <= 0;
      __delay_data_1231__delay_1230__delay_1229__delay_1228___cond_957 <= 0;
      __delay_data_1248__delay_1247__delay_1246__delay_1245___cond_964 <= 0;
      __delay_data_1265__delay_1264__delay_1263___plus_1025 <= 0;
      __delay_data_1283__delay_1282__delay_1281__delay_1280_eq_1031 <= 0;
      __delay_data_1312__delay_1311__delay_1310__delay_1309_eq_1034 <= 0;
      __delay_data_1200__delay_1199__delay_1198____variable_941 <= 0;
      __delay_data_1210__delay_1209__delay_1208___plus_1020 <= 0;
      __delay_data_1221__delay_1220__delay_1219____variable_936 <= 0;
      __delay_data_1232__delay_1231__delay_1230__delay_1229___cond_957 <= 0;
      __delay_data_1249__delay_1248__delay_1247__delay_1246___cond_964 <= 0;
      __delay_data_1266__delay_1265__delay_1264___plus_1025 <= 0;
      __delay_data_1284__delay_1283__delay_1282__delay_1281___eq_1031 <= 0;
      __delay_data_1313__delay_1312__delay_1311__delay_1310___eq_1034 <= 0;
      __delay_data_1201__delay_1200__delay_1199____variable_941 <= 0;
      __delay_data_1211__delay_1210__delay_1209___plus_1020 <= 0;
      __delay_data_1222__delay_1221__delay_1220____variable_936 <= 0;
      __delay_data_1233__delay_1232__delay_1231__delay_1230___cond_957 <= 0;
      __delay_data_1250__delay_1249__delay_1248__delay_1247___cond_964 <= 0;
      __delay_data_1267__delay_1266__delay_1265___plus_1025 <= 0;
      __delay_data_1285__delay_1284__delay_1283__delay_1282___eq_1031 <= 0;
      __delay_data_1314__delay_1313__delay_1312__delay_1311___eq_1034 <= 0;
      __delay_data_1202__delay_1201__delay_1200____variable_941 <= 0;
      __delay_data_1212__delay_1211__delay_1210___plus_1020 <= 0;
      __delay_data_1223__delay_1222__delay_1221____variable_936 <= 0;
      __delay_data_1234__delay_1233__delay_1232__delay_1231___cond_957 <= 0;
      __delay_data_1251__delay_1250__delay_1249__delay_1248___cond_964 <= 0;
      __delay_data_1268__delay_1267__delay_1266___plus_1025 <= 0;
      __delay_data_1286__delay_1285__delay_1284__delay_1283___eq_1031 <= 0;
      __delay_data_1315__delay_1314__delay_1313__delay_1312___eq_1034 <= 0;
      __delay_data_1203__delay_1202__delay_1201____variable_941 <= 0;
      __delay_data_1213__delay_1212__delay_1211___plus_1020 <= 0;
      __delay_data_1224__delay_1223__delay_1222____variable_936 <= 0;
      __delay_data_1235__delay_1234__delay_1233__delay_1232___cond_957 <= 0;
      __delay_data_1252__delay_1251__delay_1250__delay_1249___cond_964 <= 0;
      __delay_data_1269__delay_1268__delay_1267___plus_1025 <= 0;
      __delay_data_1287__delay_1286__delay_1285__delay_1284___eq_1031 <= 0;
      __delay_data_1316__delay_1315__delay_1314__delay_1313___eq_1034 <= 0;
      __delay_data_1204__delay_1203__delay_1202____variable_941 <= 0;
      __delay_data_1214__delay_1213__delay_1212___plus_1020 <= 0;
      __delay_data_1225__delay_1224__delay_1223____variable_936 <= 0;
      __delay_data_1236__delay_1235__delay_1234__delay_1233___cond_957 <= 0;
      __delay_data_1253__delay_1252__delay_1251__delay_1250___cond_964 <= 0;
      __delay_data_1270__delay_1269__delay_1268___plus_1025 <= 0;
      __delay_data_1288__delay_1287__delay_1286__delay_1285___eq_1031 <= 0;
      __delay_data_1317__delay_1316__delay_1315__delay_1314___eq_1034 <= 0;
      __delay_data_1205__delay_1204__delay_1203____variable_941 <= 0;
      __delay_data_1215__delay_1214__delay_1213___plus_1020 <= 0;
      __delay_data_1226__delay_1225__delay_1224____variable_936 <= 0;
      __delay_data_1237__delay_1236__delay_1235__delay_1234___cond_957 <= 0;
      __delay_data_1254__delay_1253__delay_1252__delay_1251___cond_964 <= 0;
      __delay_data_1271__delay_1270__delay_1269___plus_1025 <= 0;
      __delay_data_1289__delay_1288__delay_1287__delay_1286___eq_1031 <= 0;
      __delay_data_1318__delay_1317__delay_1316__delay_1315___eq_1034 <= 0;
      __delay_data_1238__delay_1237__delay_1236__delay_1235___cond_957 <= 0;
      __delay_data_1255__delay_1254__delay_1253__delay_1252___cond_964 <= 0;
      __delay_data_1272__delay_1271__delay_1270___plus_1025 <= 0;
      __delay_data_1290__delay_1289__delay_1288__delay_1287___eq_1031 <= 0;
      __delay_data_1319__delay_1318__delay_1317__delay_1316___eq_1034 <= 0;
      __delay_data_1239__delay_1238__delay_1237__delay_1236___cond_957 <= 0;
      __delay_data_1256__delay_1255__delay_1254__delay_1253___cond_964 <= 0;
      __delay_data_1273__delay_1272__delay_1271___plus_1025 <= 0;
      __delay_data_1291__delay_1290__delay_1289__delay_1288___eq_1031 <= 0;
      __delay_data_1320__delay_1319__delay_1318__delay_1317___eq_1034 <= 0;
      __delay_data_1240__delay_1239__delay_1238__delay_1237___cond_957 <= 0;
      __delay_data_1257__delay_1256__delay_1255__delay_1254___cond_964 <= 0;
      __delay_data_1274__delay_1273__delay_1272___plus_1025 <= 0;
      __delay_data_1292__delay_1291__delay_1290__delay_1289___eq_1031 <= 0;
      __delay_data_1321__delay_1320__delay_1319__delay_1318___eq_1034 <= 0;
      __delay_data_1241__delay_1240__delay_1239__delay_1238___cond_957 <= 0;
      __delay_data_1258__delay_1257__delay_1256__delay_1255___cond_964 <= 0;
      __delay_data_1275__delay_1274__delay_1273___plus_1025 <= 0;
      __delay_data_1293__delay_1292__delay_1291__delay_1290___eq_1031 <= 0;
      __delay_data_1322__delay_1321__delay_1320__delay_1319___eq_1034 <= 0;
      __delay_data_1242__delay_1241__delay_1240__delay_1239___cond_957 <= 0;
      __delay_data_1259__delay_1258__delay_1257__delay_1256___cond_964 <= 0;
      __delay_data_1276__delay_1275__delay_1274___plus_1025 <= 0;
      __delay_data_1294__delay_1293__delay_1292__delay_1291___eq_1031 <= 0;
      __delay_data_1323__delay_1322__delay_1321__delay_1320___eq_1034 <= 0;
      __delay_data_1243__delay_1242__delay_1241__delay_1240___cond_957 <= 0;
      __delay_data_1260__delay_1259__delay_1258__delay_1257___cond_964 <= 0;
      __delay_data_1277__delay_1276__delay_1275___plus_1025 <= 0;
      __delay_data_1295__delay_1294__delay_1293__delay_1292___eq_1031 <= 0;
      __delay_data_1324__delay_1323__delay_1322__delay_1321___eq_1034 <= 0;
      _plus_data_1023 <= 0;
      __delay_data_1261__delay_1260__delay_1259__delay_1258___cond_964 <= 0;
      __delay_data_1278__delay_1277__delay_1276___plus_1025 <= 0;
      __delay_data_1296__delay_1295__delay_1294__delay_1293___eq_1031 <= 0;
      __delay_data_1325__delay_1324__delay_1323__delay_1322___eq_1034 <= 0;
      __delay_data_1337__substreamoutput_1022 <= 0;
      __delay_data_1297__delay_1296__delay_1295__delay_1294___eq_1031 <= 0;
      __delay_data_1326__delay_1325__delay_1324__delay_1323___eq_1034 <= 0;
      __delay_data_1338__delay_1337__substreamoutput_1022 <= 0;
      __delay_data_1298__delay_1297__delay_1296__delay_1295___eq_1031 <= 0;
      __delay_data_1327__delay_1326__delay_1325__delay_1324___eq_1034 <= 0;
      __delay_data_1339__delay_1338____substreamoutput_1022 <= 0;
      __delay_data_1299__delay_1298__delay_1297__delay_1296___eq_1031 <= 0;
      __delay_data_1328__delay_1327__delay_1326__delay_1325___eq_1034 <= 0;
      __delay_data_1340__delay_1339____substreamoutput_1022 <= 0;
      __delay_data_1300__delay_1299__delay_1298__delay_1297___eq_1031 <= 0;
      __delay_data_1329__delay_1328__delay_1327__delay_1326___eq_1034 <= 0;
      __delay_data_1341__delay_1340____substreamoutput_1022 <= 0;
      __delay_data_1301__delay_1300__delay_1299__delay_1298___eq_1031 <= 0;
      __delay_data_1330__delay_1329__delay_1328__delay_1327___eq_1034 <= 0;
      __delay_data_1342__delay_1341____substreamoutput_1022 <= 0;
      __delay_data_1302__delay_1301__delay_1300__delay_1299___eq_1031 <= 0;
      __delay_data_1331__delay_1330__delay_1329__delay_1328___eq_1034 <= 0;
      __delay_data_1343__delay_1342____substreamoutput_1022 <= 0;
      __delay_data_1303__delay_1302__delay_1301__delay_1300___eq_1031 <= 0;
      __delay_data_1332__delay_1331__delay_1330__delay_1329___eq_1034 <= 0;
      __delay_data_1344__delay_1343____substreamoutput_1022 <= 0;
      __delay_data_1304__delay_1303__delay_1302__delay_1301___eq_1031 <= 0;
      __delay_data_1333__delay_1332__delay_1331__delay_1330___eq_1034 <= 0;
      __delay_data_1345__delay_1344____substreamoutput_1022 <= 0;
      __delay_data_1305__delay_1304__delay_1303__delay_1302___eq_1031 <= 0;
      __delay_data_1334__delay_1333__delay_1332__delay_1331___eq_1034 <= 0;
      __delay_data_1346__delay_1345____substreamoutput_1022 <= 0;
      _greaterthan_data_1028 <= 0;
      __delay_data_1279__substreamoutput_1026 <= 0;
      __delay_data_1306__delay_1305__delay_1304__delay_1303___eq_1031 <= 0;
      __delay_data_1335__delay_1334__delay_1333__delay_1332___eq_1034 <= 0;
      __delay_data_1347__delay_1346____substreamoutput_1022 <= 0;
      _cond_data_1030 <= 0;
      __delay_data_1307__delay_1306__delay_1305__delay_1304___eq_1031 <= 0;
      __delay_data_1308__delay_1279__substreamoutput_1026 <= 0;
      __delay_data_1336__delay_1335__delay_1334__delay_1333___eq_1034 <= 0;
      __delay_data_1348__delay_1347____substreamoutput_1022 <= 0;
      _stream_matmul_55_parameter_0_next_parameter_data <= 0;
      __variable_wdata_936 <= 0;
      _stream_matmul_55_parameter_1_next_parameter_data <= 0;
      __variable_wdata_937 <= 0;
      _stream_matmul_55_parameter_2_next_parameter_data <= 0;
      __variable_wdata_938 <= 0;
      _stream_matmul_55_parameter_3_next_parameter_data <= 0;
      __variable_wdata_939 <= 0;
      _stream_matmul_55_parameter_4_next_parameter_data <= 0;
      __variable_wdata_940 <= 0;
      _stream_matmul_55_parameter_6_next_parameter_data <= 0;
      __variable_wdata_951 <= 0;
      _stream_matmul_55_source_7_source_mode <= 5'b0;
      _stream_matmul_55_source_7_source_offset <= 0;
      _source_stream_matmul_55_source_7_pat_size_0 <= 0;
      _source_stream_matmul_55_source_7_pat_stride_0 <= 0;
      _source_stream_matmul_55_source_7_pat_size_1 <= 0;
      _source_stream_matmul_55_source_7_pat_stride_1 <= 0;
      _source_stream_matmul_55_source_7_pat_size_2 <= 0;
      _source_stream_matmul_55_source_7_pat_stride_2 <= 0;
      _source_stream_matmul_55_source_7_pat_size_3 <= 0;
      _source_stream_matmul_55_source_7_pat_stride_3 <= 0;
      _stream_matmul_55_source_7_source_sel <= 0;
      _stream_matmul_55_source_7_source_offset_buf <= 0;
      _source_stream_matmul_55_source_7_pat_cur_offset_0 <= 0;
      _source_stream_matmul_55_source_7_pat_cur_offset_1 <= 0;
      _source_stream_matmul_55_source_7_pat_cur_offset_2 <= 0;
      _source_stream_matmul_55_source_7_pat_cur_offset_3 <= 0;
      _source_stream_matmul_55_source_7_pat_count_0 <= 0;
      _source_stream_matmul_55_source_7_pat_count_1 <= 0;
      _source_stream_matmul_55_source_7_pat_count_2 <= 0;
      _source_stream_matmul_55_source_7_pat_count_3 <= 0;
      _source_stream_matmul_55_source_7_pat_size_buf_0 <= 0;
      _source_stream_matmul_55_source_7_pat_size_buf_1 <= 0;
      _source_stream_matmul_55_source_7_pat_size_buf_2 <= 0;
      _source_stream_matmul_55_source_7_pat_size_buf_3 <= 0;
      _source_stream_matmul_55_source_7_pat_stride_buf_0 <= 0;
      _source_stream_matmul_55_source_7_pat_stride_buf_1 <= 0;
      _source_stream_matmul_55_source_7_pat_stride_buf_2 <= 0;
      _source_stream_matmul_55_source_7_pat_stride_buf_3 <= 0;
      __variable_wdata_952 <= 0;
      _stream_matmul_55_source_7_source_ram_raddr <= 0;
      _stream_matmul_55_parameter_8_next_parameter_data <= 0;
      __variable_wdata_958 <= 0;
      _stream_matmul_55_source_9_source_mode <= 5'b0;
      _stream_matmul_55_source_9_source_offset <= 0;
      _source_stream_matmul_55_source_9_pat_size_0 <= 0;
      _source_stream_matmul_55_source_9_pat_stride_0 <= 0;
      _source_stream_matmul_55_source_9_pat_size_1 <= 0;
      _source_stream_matmul_55_source_9_pat_stride_1 <= 0;
      _source_stream_matmul_55_source_9_pat_size_2 <= 0;
      _source_stream_matmul_55_source_9_pat_stride_2 <= 0;
      _source_stream_matmul_55_source_9_pat_size_3 <= 0;
      _source_stream_matmul_55_source_9_pat_stride_3 <= 0;
      _stream_matmul_55_source_9_source_sel <= 0;
      _stream_matmul_55_source_9_source_offset_buf <= 0;
      _source_stream_matmul_55_source_9_pat_cur_offset_0 <= 0;
      _source_stream_matmul_55_source_9_pat_cur_offset_1 <= 0;
      _source_stream_matmul_55_source_9_pat_cur_offset_2 <= 0;
      _source_stream_matmul_55_source_9_pat_cur_offset_3 <= 0;
      _source_stream_matmul_55_source_9_pat_count_0 <= 0;
      _source_stream_matmul_55_source_9_pat_count_1 <= 0;
      _source_stream_matmul_55_source_9_pat_count_2 <= 0;
      _source_stream_matmul_55_source_9_pat_count_3 <= 0;
      _source_stream_matmul_55_source_9_pat_size_buf_0 <= 0;
      _source_stream_matmul_55_source_9_pat_size_buf_1 <= 0;
      _source_stream_matmul_55_source_9_pat_size_buf_2 <= 0;
      _source_stream_matmul_55_source_9_pat_size_buf_3 <= 0;
      _source_stream_matmul_55_source_9_pat_stride_buf_0 <= 0;
      _source_stream_matmul_55_source_9_pat_stride_buf_1 <= 0;
      _source_stream_matmul_55_source_9_pat_stride_buf_2 <= 0;
      _source_stream_matmul_55_source_9_pat_stride_buf_3 <= 0;
      __variable_wdata_959 <= 0;
      _stream_matmul_55_source_9_source_ram_raddr <= 0;
      _stream_matmul_55_parameter_10_next_parameter_data <= 0;
      __variable_wdata_965 <= 0;
      _stream_matmul_55_source_11_source_mode <= 5'b0;
      _stream_matmul_55_source_11_source_empty_data <= 0;
      __variable_wdata_966 <= 0;
      _stream_matmul_55_parameter_12_next_parameter_data <= 0;
      __variable_wdata_972 <= 0;
      _stream_matmul_55_source_13_source_mode <= 5'b0;
      _stream_matmul_55_source_13_source_empty_data <= 0;
      __variable_wdata_973 <= 0;
      _stream_matmul_55_parameter_14_next_parameter_data <= 0;
      __variable_wdata_979 <= 0;
      _stream_matmul_55_source_15_source_mode <= 5'b0;
      _stream_matmul_55_source_15_source_empty_data <= 0;
      __variable_wdata_980 <= 0;
      _stream_matmul_55_parameter_16_next_parameter_data <= 0;
      __variable_wdata_986 <= 0;
      _stream_matmul_55_parameter_17_next_parameter_data <= 0;
      __variable_wdata_987 <= 0;
      _stream_matmul_55_parameter_18_next_parameter_data <= 0;
      __variable_wdata_988 <= 0;
      _stream_matmul_55_parameter_19_next_parameter_data <= 0;
      __variable_wdata_989 <= 0;
      _stream_matmul_55_source_20_source_mode <= 5'b0;
      _stream_matmul_55_source_20_source_offset <= 0;
      _source_stream_matmul_55_source_20_pat_size_0 <= 0;
      _source_stream_matmul_55_source_20_pat_stride_0 <= 0;
      _source_stream_matmul_55_source_20_pat_size_1 <= 0;
      _source_stream_matmul_55_source_20_pat_stride_1 <= 0;
      _source_stream_matmul_55_source_20_pat_size_2 <= 0;
      _source_stream_matmul_55_source_20_pat_stride_2 <= 0;
      _source_stream_matmul_55_source_20_pat_size_3 <= 0;
      _source_stream_matmul_55_source_20_pat_stride_3 <= 0;
      _stream_matmul_55_source_20_source_sel <= 0;
      _stream_matmul_55_source_20_source_offset_buf <= 0;
      _source_stream_matmul_55_source_20_pat_cur_offset_0 <= 0;
      _source_stream_matmul_55_source_20_pat_cur_offset_1 <= 0;
      _source_stream_matmul_55_source_20_pat_cur_offset_2 <= 0;
      _source_stream_matmul_55_source_20_pat_cur_offset_3 <= 0;
      _source_stream_matmul_55_source_20_pat_count_0 <= 0;
      _source_stream_matmul_55_source_20_pat_count_1 <= 0;
      _source_stream_matmul_55_source_20_pat_count_2 <= 0;
      _source_stream_matmul_55_source_20_pat_count_3 <= 0;
      _source_stream_matmul_55_source_20_pat_size_buf_0 <= 0;
      _source_stream_matmul_55_source_20_pat_size_buf_1 <= 0;
      _source_stream_matmul_55_source_20_pat_size_buf_2 <= 0;
      _source_stream_matmul_55_source_20_pat_size_buf_3 <= 0;
      _source_stream_matmul_55_source_20_pat_stride_buf_0 <= 0;
      _source_stream_matmul_55_source_20_pat_stride_buf_1 <= 0;
      _source_stream_matmul_55_source_20_pat_stride_buf_2 <= 0;
      _source_stream_matmul_55_source_20_pat_stride_buf_3 <= 0;
      __variable_wdata_990 <= 0;
      _stream_matmul_55_source_20_source_ram_raddr <= 0;
      _stream_matmul_55_source_21_source_mode <= 5'b0;
      _stream_matmul_55_source_21_source_offset <= 0;
      _source_stream_matmul_55_source_21_pat_size_0 <= 0;
      _source_stream_matmul_55_source_21_pat_stride_0 <= 0;
      _source_stream_matmul_55_source_21_pat_size_1 <= 0;
      _source_stream_matmul_55_source_21_pat_stride_1 <= 0;
      _source_stream_matmul_55_source_21_pat_size_2 <= 0;
      _source_stream_matmul_55_source_21_pat_stride_2 <= 0;
      _source_stream_matmul_55_source_21_pat_size_3 <= 0;
      _source_stream_matmul_55_source_21_pat_stride_3 <= 0;
      _stream_matmul_55_source_21_source_sel <= 0;
      _stream_matmul_55_source_21_source_offset_buf <= 0;
      _source_stream_matmul_55_source_21_pat_cur_offset_0 <= 0;
      _source_stream_matmul_55_source_21_pat_cur_offset_1 <= 0;
      _source_stream_matmul_55_source_21_pat_cur_offset_2 <= 0;
      _source_stream_matmul_55_source_21_pat_cur_offset_3 <= 0;
      _source_stream_matmul_55_source_21_pat_count_0 <= 0;
      _source_stream_matmul_55_source_21_pat_count_1 <= 0;
      _source_stream_matmul_55_source_21_pat_count_2 <= 0;
      _source_stream_matmul_55_source_21_pat_count_3 <= 0;
      _source_stream_matmul_55_source_21_pat_size_buf_0 <= 0;
      _source_stream_matmul_55_source_21_pat_size_buf_1 <= 0;
      _source_stream_matmul_55_source_21_pat_size_buf_2 <= 0;
      _source_stream_matmul_55_source_21_pat_size_buf_3 <= 0;
      _source_stream_matmul_55_source_21_pat_stride_buf_0 <= 0;
      _source_stream_matmul_55_source_21_pat_stride_buf_1 <= 0;
      _source_stream_matmul_55_source_21_pat_stride_buf_2 <= 0;
      _source_stream_matmul_55_source_21_pat_stride_buf_3 <= 0;
      __variable_wdata_1004 <= 0;
      _stream_matmul_55_source_21_source_ram_raddr <= 0;
      _tmp_1716 <= 0;
      _tmp_1717 <= 0;
      _tmp_1718 <= 0;
      _tmp_1719 <= 0;
      _tmp_1720 <= 0;
      _tmp_1721 <= 0;
      _tmp_1722 <= 0;
      _tmp_1723 <= 0;
      _tmp_1724 <= 0;
      _tmp_1725 <= 0;
      _tmp_1726 <= 0;
      _tmp_1727 <= 0;
      _tmp_1728 <= 0;
      _tmp_1729 <= 0;
      _tmp_1730 <= 0;
      _tmp_1731 <= 0;
      _tmp_1732 <= 0;
      _tmp_1733 <= 0;
      _tmp_1734 <= 0;
      _tmp_1735 <= 0;
      _tmp_1736 <= 0;
      _tmp_1737 <= 0;
      _tmp_1738 <= 0;
      _tmp_1739 <= 0;
      _tmp_1740 <= 0;
      _tmp_1741 <= 0;
      _tmp_1742 <= 0;
      _tmp_1743 <= 0;
      _tmp_1744 <= 0;
      _tmp_1745 <= 0;
      _tmp_1746 <= 0;
      _tmp_1749 <= 0;
      _tmp_1750 <= 0;
      _tmp_1751 <= 0;
      _tmp_1752 <= 0;
      _tmp_1753 <= 0;
      _tmp_1754 <= 0;
      _tmp_1755 <= 0;
      _tmp_1756 <= 0;
      _tmp_1757 <= 0;
      _tmp_1758 <= 0;
      _tmp_1759 <= 0;
      _tmp_1760 <= 0;
      _tmp_1761 <= 0;
      _tmp_1762 <= 0;
      _tmp_1763 <= 0;
      _tmp_1764 <= 0;
      _tmp_1765 <= 0;
      _tmp_1766 <= 0;
      _tmp_1767 <= 0;
      _tmp_1768 <= 0;
      _tmp_1769 <= 0;
      _tmp_1770 <= 0;
      _tmp_1771 <= 0;
      _tmp_1772 <= 0;
      _tmp_1773 <= 0;
      _tmp_1774 <= 0;
      _tmp_1775 <= 0;
      _tmp_1776 <= 0;
      _tmp_1777 <= 0;
      _tmp_1778 <= 0;
      _tmp_1779 <= 0;
      _tmp_1780 <= 0;
      _tmp_1781 <= 0;
      _tmp_1782 <= 0;
      _tmp_1783 <= 0;
      _tmp_1784 <= 0;
      _tmp_1785 <= 0;
      _tmp_1786 <= 0;
      _tmp_1787 <= 0;
      _tmp_1788 <= 0;
      _tmp_1789 <= 0;
      _tmp_1790 <= 0;
      _tmp_1791 <= 0;
      _tmp_1792 <= 0;
      _tmp_1793 <= 0;
      _tmp_1794 <= 0;
      _tmp_1795 <= 0;
      _tmp_1796 <= 0;
      _tmp_1797 <= 0;
      _tmp_1798 <= 0;
      _tmp_1799 <= 0;
      _tmp_1800 <= 0;
      _tmp_1801 <= 0;
      _tmp_1802 <= 0;
      _tmp_1803 <= 0;
      _tmp_1804 <= 0;
      _tmp_1805 <= 0;
      _tmp_1806 <= 0;
      _tmp_1807 <= 0;
      _tmp_1808 <= 0;
      _tmp_1809 <= 0;
      _tmp_1810 <= 0;
      _stream_matmul_55_sink_26_sink_mode <= 5'b0;
      _stream_matmul_55_sink_26_sink_offset <= 0;
      _stream_matmul_55_sink_26_sink_size <= 0;
      _stream_matmul_55_sink_26_sink_stride <= 0;
      _stream_matmul_55_sink_26_sink_sel <= 0;
      _stream_matmul_55_sink_26_sink_offset_buf <= 0;
      _stream_matmul_55_sink_26_sink_size_buf <= 0;
      _stream_matmul_55_sink_26_sink_stride_buf <= 0;
      _stream_matmul_55_sink_26_sink_waddr <= 0;
      _stream_matmul_55_sink_26_sink_count <= 0;
      _stream_matmul_55_sink_26_sink_wdata <= 0;
      _tmp_1823 <= 0;
      _tmp_1824 <= 0;
      _tmp_1825 <= 0;
      _tmp_1826 <= 0;
      _tmp_1827 <= 0;
      _tmp_1828 <= 0;
      __variable_wdata_941 <= 0;
      _tmp_1829 <= 0;
      _tmp_1830 <= 0;
      _tmp_1831 <= 0;
      _tmp_1832 <= 0;
      _tmp_1835 <= 0;
      _tmp_1838 <= 0;
      _tmp_1839 <= 0;
      _tmp_1840 <= 0;
      _tmp_1841 <= 0;
      _tmp_1842 <= 0;
      _tmp_1843 <= 0;
      _tmp_1844 <= 0;
      _tmp_1845 <= 0;
      _tmp_1846 <= 0;
      _tmp_1847 <= 0;
      _tmp_1848 <= 0;
      _tmp_1849 <= 0;
      _tmp_1850 <= 0;
      _tmp_1851 <= 0;
      _tmp_1852 <= 0;
      _tmp_1853 <= 0;
      _tmp_1854 <= 0;
      _tmp_1855 <= 0;
      _tmp_1856 <= 0;
      _tmp_1857 <= 0;
      _tmp_1858 <= 0;
      _tmp_1859 <= 0;
      _tmp_1860 <= 0;
      _tmp_1861 <= 0;
      _tmp_1862 <= 0;
      _tmp_1863 <= 0;
      _tmp_1864 <= 0;
      _tmp_1865 <= 0;
      _tmp_1866 <= 0;
      _tmp_1867 <= 0;
      _tmp_1868 <= 0;
      _tmp_1869 <= 0;
      _tmp_1870 <= 0;
      _tmp_1871 <= 0;
      _tmp_1872 <= 0;
      _tmp_1873 <= 0;
      _tmp_1874 <= 0;
      _tmp_1875 <= 0;
      _tmp_1876 <= 0;
      _tmp_1877 <= 0;
      _tmp_1878 <= 0;
      _tmp_1879 <= 0;
      _tmp_1880 <= 0;
      _tmp_1881 <= 0;
      _tmp_1882 <= 0;
      _tmp_1883 <= 0;
      _tmp_1884 <= 0;
      _tmp_1885 <= 0;
      _tmp_1886 <= 0;
      _tmp_1887 <= 0;
      _tmp_1888 <= 0;
      _tmp_1889 <= 0;
      _tmp_1890 <= 0;
      _tmp_1891 <= 0;
      _tmp_1892 <= 0;
      _tmp_1893 <= 0;
      _tmp_1894 <= 0;
      _tmp_1895 <= 0;
      _tmp_1896 <= 0;
      _tmp_1897 <= 0;
      _tmp_1898 <= 0;
      _tmp_1899 <= 0;
      _tmp_1900 <= 0;
      _tmp_1901 <= 0;
      _tmp_1902 <= 0;
      _tmp_1903 <= 0;
      _tmp_1904 <= 0;
      _tmp_1905 <= 0;
      _tmp_1906 <= 0;
      _tmp_1907 <= 0;
      _tmp_1908 <= 0;
      _tmp_1909 <= 0;
      _tmp_1910 <= 0;
      _tmp_1911 <= 0;
      _tmp_1912 <= 0;
      _tmp_1913 <= 0;
      _tmp_1914 <= 0;
      _tmp_1915 <= 0;
      _tmp_1916 <= 0;
      _tmp_1917 <= 0;
      _tmp_1918 <= 0;
      _tmp_1919 <= 0;
      _tmp_1920 <= 0;
      _tmp_1921 <= 0;
      _tmp_1922 <= 0;
      _tmp_1923 <= 0;
      _tmp_1924 <= 0;
      _tmp_1925 <= 0;
      _tmp_1926 <= 0;
      _tmp_1927 <= 0;
      _tmp_1928 <= 0;
      _tmp_1929 <= 0;
      _tmp_1930 <= 0;
      _tmp_1931 <= 0;
      _tmp_1932 <= 0;
      _stream_matmul_55_busy_reg <= 0;
    end else begin
      if(_stream_matmul_55_stream_oready) begin
        _stream_matmul_55_source_7_source_ram_renable <= 0;
        _stream_matmul_55_source_7_source_fifo_deq <= 0;
      end 
      _stream_matmul_55_source_7_idle <= _stream_matmul_55_source_7_idle;
      if(_stream_matmul_55_stream_oready) begin
        _stream_matmul_55_source_9_source_ram_renable <= 0;
        _stream_matmul_55_source_9_source_fifo_deq <= 0;
      end 
      _stream_matmul_55_source_9_idle <= _stream_matmul_55_source_9_idle;
      if(_stream_matmul_55_stream_oready) begin
        _stream_matmul_55_source_11_source_ram_renable <= 0;
        _stream_matmul_55_source_11_source_fifo_deq <= 0;
      end 
      _stream_matmul_55_source_11_idle <= _stream_matmul_55_source_11_idle;
      if(_stream_matmul_55_stream_oready) begin
        _stream_matmul_55_source_13_source_ram_renable <= 0;
        _stream_matmul_55_source_13_source_fifo_deq <= 0;
      end 
      _stream_matmul_55_source_13_idle <= _stream_matmul_55_source_13_idle;
      if(_stream_matmul_55_stream_oready) begin
        _stream_matmul_55_source_15_source_ram_renable <= 0;
        _stream_matmul_55_source_15_source_fifo_deq <= 0;
      end 
      _stream_matmul_55_source_15_idle <= _stream_matmul_55_source_15_idle;
      if(_stream_matmul_55_stream_oready) begin
        _stream_matmul_55_source_20_source_ram_renable <= 0;
        _stream_matmul_55_source_20_source_fifo_deq <= 0;
      end 
      _stream_matmul_55_source_20_idle <= _stream_matmul_55_source_20_idle;
      if(_stream_matmul_55_stream_oready) begin
        _stream_matmul_55_source_21_source_ram_renable <= 0;
        _stream_matmul_55_source_21_source_fifo_deq <= 0;
      end 
      _stream_matmul_55_source_21_idle <= _stream_matmul_55_source_21_idle;
      if(_stream_matmul_55_stream_oready) begin
        _stream_matmul_55_sink_26_sink_wenable <= 0;
        _stream_matmul_55_sink_26_sink_fifo_enq <= 0;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _stream_matmul_55_sink_27_sink_wenable <= 0;
        _stream_matmul_55_sink_27_sink_fifo_enq <= 0;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __stream_matmul_55_stream_ivalid_1 <= _stream_matmul_55_stream_ivalid;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __stream_matmul_55_stream_ivalid_2 <= __stream_matmul_55_stream_ivalid_1;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __stream_matmul_55_stream_ivalid_3 <= __stream_matmul_55_stream_ivalid_2;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __stream_matmul_55_stream_ivalid_4 <= __stream_matmul_55_stream_ivalid_3;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __stream_matmul_55_stream_ivalid_5 <= __stream_matmul_55_stream_ivalid_4;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __stream_matmul_55_stream_ivalid_6 <= __stream_matmul_55_stream_ivalid_5;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __stream_matmul_55_stream_ivalid_7 <= __stream_matmul_55_stream_ivalid_6;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __stream_matmul_55_stream_ivalid_8 <= __stream_matmul_55_stream_ivalid_7;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __stream_matmul_55_stream_ivalid_9 <= __stream_matmul_55_stream_ivalid_8;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __stream_matmul_55_stream_ivalid_10 <= __stream_matmul_55_stream_ivalid_9;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __stream_matmul_55_stream_ivalid_11 <= __stream_matmul_55_stream_ivalid_10;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __stream_matmul_55_stream_ivalid_12 <= __stream_matmul_55_stream_ivalid_11;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __stream_matmul_55_stream_ivalid_13 <= __stream_matmul_55_stream_ivalid_12;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __stream_matmul_55_stream_ivalid_14 <= __stream_matmul_55_stream_ivalid_13;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __stream_matmul_55_stream_ivalid_15 <= __stream_matmul_55_stream_ivalid_14;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __stream_matmul_55_stream_ivalid_16 <= __stream_matmul_55_stream_ivalid_15;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __stream_matmul_55_stream_ivalid_17 <= __stream_matmul_55_stream_ivalid_16;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __stream_matmul_55_stream_ivalid_18 <= __stream_matmul_55_stream_ivalid_17;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __stream_matmul_55_stream_ivalid_19 <= __stream_matmul_55_stream_ivalid_18;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __stream_matmul_55_stream_ivalid_20 <= __stream_matmul_55_stream_ivalid_19;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __stream_matmul_55_stream_ivalid_21 <= __stream_matmul_55_stream_ivalid_20;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __stream_matmul_55_stream_ivalid_22 <= __stream_matmul_55_stream_ivalid_21;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __stream_matmul_55_stream_ivalid_23 <= __stream_matmul_55_stream_ivalid_22;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __stream_matmul_55_stream_ivalid_24 <= __stream_matmul_55_stream_ivalid_23;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __stream_matmul_55_stream_ivalid_25 <= __stream_matmul_55_stream_ivalid_24;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __stream_matmul_55_stream_ivalid_26 <= __stream_matmul_55_stream_ivalid_25;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __stream_matmul_55_stream_ivalid_27 <= __stream_matmul_55_stream_ivalid_26;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __stream_matmul_55_stream_ivalid_28 <= __stream_matmul_55_stream_ivalid_27;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __stream_matmul_55_stream_ivalid_29 <= __stream_matmul_55_stream_ivalid_28;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _eq_data_991 <= stream_matmul_55_parameter_1_data == 1'sd0;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _eq_data_995 <= stream_matmul_55_parameter_2_data == 1'sd0;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _plus_data_1015 <= _cond_data_971 + stream_matmul_55_parameter_16_data;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _plus_data_1020 <= _cond_data_978 + stream_matmul_55_parameter_17_data;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _plus_data_1025 <= _cond_data_985 + stream_matmul_55_parameter_18_data;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _eq_data_1031 <= stream_matmul_55_parameter_19_data == 1'sd0;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _eq_data_1034 <= stream_matmul_55_parameter_19_data == 2'sd1;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1192__variable_990 <= stream_matmul_55_source_20_data;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1193_pointer_1010 <= _pointer_data_1010;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1194_reinterpretcast_1009 <= _reinterpretcast_data_1009;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1195__variable_941 <= stream_matmul_55__reduce_reset_data;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1216__variable_936 <= stream_matmul_55_parameter_0_data;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1227_cond_957 <= _cond_data_957;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1244_cond_964 <= _cond_data_964;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1196__delay_1195__variable_941 <= __delay_data_1195__variable_941;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1206_plus_1020 <= _plus_data_1020;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1217__delay_1216__variable_936 <= __delay_data_1216__variable_936;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1228__delay_1227_cond_957 <= __delay_data_1227_cond_957;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1245__delay_1244_cond_964 <= __delay_data_1244_cond_964;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1262_plus_1025 <= _plus_data_1025;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1280_eq_1031 <= _eq_data_1031;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1309_eq_1034 <= _eq_data_1034;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1197__delay_1196__delay_1195__variable_941 <= __delay_data_1196__delay_1195__variable_941;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1207__delay_1206_plus_1020 <= __delay_data_1206_plus_1020;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1218__delay_1217__delay_1216__variable_936 <= __delay_data_1217__delay_1216__variable_936;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1229__delay_1228__delay_1227_cond_957 <= __delay_data_1228__delay_1227_cond_957;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1246__delay_1245__delay_1244_cond_964 <= __delay_data_1245__delay_1244_cond_964;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1263__delay_1262_plus_1025 <= __delay_data_1262_plus_1025;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1281__delay_1280_eq_1031 <= __delay_data_1280_eq_1031;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1310__delay_1309_eq_1034 <= __delay_data_1309_eq_1034;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1198__delay_1197__delay_1196____variable_941 <= __delay_data_1197__delay_1196__delay_1195__variable_941;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1208__delay_1207__delay_1206_plus_1020 <= __delay_data_1207__delay_1206_plus_1020;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1219__delay_1218__delay_1217____variable_936 <= __delay_data_1218__delay_1217__delay_1216__variable_936;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1230__delay_1229__delay_1228__delay_1227_cond_957 <= __delay_data_1229__delay_1228__delay_1227_cond_957;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1247__delay_1246__delay_1245__delay_1244_cond_964 <= __delay_data_1246__delay_1245__delay_1244_cond_964;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1264__delay_1263__delay_1262_plus_1025 <= __delay_data_1263__delay_1262_plus_1025;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1282__delay_1281__delay_1280_eq_1031 <= __delay_data_1281__delay_1280_eq_1031;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1311__delay_1310__delay_1309_eq_1034 <= __delay_data_1310__delay_1309_eq_1034;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1199__delay_1198__delay_1197____variable_941 <= __delay_data_1198__delay_1197__delay_1196____variable_941;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1209__delay_1208__delay_1207___plus_1020 <= __delay_data_1208__delay_1207__delay_1206_plus_1020;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1220__delay_1219__delay_1218____variable_936 <= __delay_data_1219__delay_1218__delay_1217____variable_936;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1231__delay_1230__delay_1229__delay_1228___cond_957 <= __delay_data_1230__delay_1229__delay_1228__delay_1227_cond_957;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1248__delay_1247__delay_1246__delay_1245___cond_964 <= __delay_data_1247__delay_1246__delay_1245__delay_1244_cond_964;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1265__delay_1264__delay_1263___plus_1025 <= __delay_data_1264__delay_1263__delay_1262_plus_1025;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1283__delay_1282__delay_1281__delay_1280_eq_1031 <= __delay_data_1282__delay_1281__delay_1280_eq_1031;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1312__delay_1311__delay_1310__delay_1309_eq_1034 <= __delay_data_1311__delay_1310__delay_1309_eq_1034;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1200__delay_1199__delay_1198____variable_941 <= __delay_data_1199__delay_1198__delay_1197____variable_941;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1210__delay_1209__delay_1208___plus_1020 <= __delay_data_1209__delay_1208__delay_1207___plus_1020;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1221__delay_1220__delay_1219____variable_936 <= __delay_data_1220__delay_1219__delay_1218____variable_936;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1232__delay_1231__delay_1230__delay_1229___cond_957 <= __delay_data_1231__delay_1230__delay_1229__delay_1228___cond_957;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1249__delay_1248__delay_1247__delay_1246___cond_964 <= __delay_data_1248__delay_1247__delay_1246__delay_1245___cond_964;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1266__delay_1265__delay_1264___plus_1025 <= __delay_data_1265__delay_1264__delay_1263___plus_1025;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1284__delay_1283__delay_1282__delay_1281___eq_1031 <= __delay_data_1283__delay_1282__delay_1281__delay_1280_eq_1031;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1313__delay_1312__delay_1311__delay_1310___eq_1034 <= __delay_data_1312__delay_1311__delay_1310__delay_1309_eq_1034;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1201__delay_1200__delay_1199____variable_941 <= __delay_data_1200__delay_1199__delay_1198____variable_941;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1211__delay_1210__delay_1209___plus_1020 <= __delay_data_1210__delay_1209__delay_1208___plus_1020;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1222__delay_1221__delay_1220____variable_936 <= __delay_data_1221__delay_1220__delay_1219____variable_936;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1233__delay_1232__delay_1231__delay_1230___cond_957 <= __delay_data_1232__delay_1231__delay_1230__delay_1229___cond_957;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1250__delay_1249__delay_1248__delay_1247___cond_964 <= __delay_data_1249__delay_1248__delay_1247__delay_1246___cond_964;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1267__delay_1266__delay_1265___plus_1025 <= __delay_data_1266__delay_1265__delay_1264___plus_1025;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1285__delay_1284__delay_1283__delay_1282___eq_1031 <= __delay_data_1284__delay_1283__delay_1282__delay_1281___eq_1031;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1314__delay_1313__delay_1312__delay_1311___eq_1034 <= __delay_data_1313__delay_1312__delay_1311__delay_1310___eq_1034;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1202__delay_1201__delay_1200____variable_941 <= __delay_data_1201__delay_1200__delay_1199____variable_941;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1212__delay_1211__delay_1210___plus_1020 <= __delay_data_1211__delay_1210__delay_1209___plus_1020;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1223__delay_1222__delay_1221____variable_936 <= __delay_data_1222__delay_1221__delay_1220____variable_936;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1234__delay_1233__delay_1232__delay_1231___cond_957 <= __delay_data_1233__delay_1232__delay_1231__delay_1230___cond_957;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1251__delay_1250__delay_1249__delay_1248___cond_964 <= __delay_data_1250__delay_1249__delay_1248__delay_1247___cond_964;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1268__delay_1267__delay_1266___plus_1025 <= __delay_data_1267__delay_1266__delay_1265___plus_1025;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1286__delay_1285__delay_1284__delay_1283___eq_1031 <= __delay_data_1285__delay_1284__delay_1283__delay_1282___eq_1031;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1315__delay_1314__delay_1313__delay_1312___eq_1034 <= __delay_data_1314__delay_1313__delay_1312__delay_1311___eq_1034;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1203__delay_1202__delay_1201____variable_941 <= __delay_data_1202__delay_1201__delay_1200____variable_941;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1213__delay_1212__delay_1211___plus_1020 <= __delay_data_1212__delay_1211__delay_1210___plus_1020;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1224__delay_1223__delay_1222____variable_936 <= __delay_data_1223__delay_1222__delay_1221____variable_936;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1235__delay_1234__delay_1233__delay_1232___cond_957 <= __delay_data_1234__delay_1233__delay_1232__delay_1231___cond_957;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1252__delay_1251__delay_1250__delay_1249___cond_964 <= __delay_data_1251__delay_1250__delay_1249__delay_1248___cond_964;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1269__delay_1268__delay_1267___plus_1025 <= __delay_data_1268__delay_1267__delay_1266___plus_1025;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1287__delay_1286__delay_1285__delay_1284___eq_1031 <= __delay_data_1286__delay_1285__delay_1284__delay_1283___eq_1031;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1316__delay_1315__delay_1314__delay_1313___eq_1034 <= __delay_data_1315__delay_1314__delay_1313__delay_1312___eq_1034;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1204__delay_1203__delay_1202____variable_941 <= __delay_data_1203__delay_1202__delay_1201____variable_941;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1214__delay_1213__delay_1212___plus_1020 <= __delay_data_1213__delay_1212__delay_1211___plus_1020;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1225__delay_1224__delay_1223____variable_936 <= __delay_data_1224__delay_1223__delay_1222____variable_936;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1236__delay_1235__delay_1234__delay_1233___cond_957 <= __delay_data_1235__delay_1234__delay_1233__delay_1232___cond_957;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1253__delay_1252__delay_1251__delay_1250___cond_964 <= __delay_data_1252__delay_1251__delay_1250__delay_1249___cond_964;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1270__delay_1269__delay_1268___plus_1025 <= __delay_data_1269__delay_1268__delay_1267___plus_1025;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1288__delay_1287__delay_1286__delay_1285___eq_1031 <= __delay_data_1287__delay_1286__delay_1285__delay_1284___eq_1031;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1317__delay_1316__delay_1315__delay_1314___eq_1034 <= __delay_data_1316__delay_1315__delay_1314__delay_1313___eq_1034;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1205__delay_1204__delay_1203____variable_941 <= __delay_data_1204__delay_1203__delay_1202____variable_941;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1215__delay_1214__delay_1213___plus_1020 <= __delay_data_1214__delay_1213__delay_1212___plus_1020;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1226__delay_1225__delay_1224____variable_936 <= __delay_data_1225__delay_1224__delay_1223____variable_936;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1237__delay_1236__delay_1235__delay_1234___cond_957 <= __delay_data_1236__delay_1235__delay_1234__delay_1233___cond_957;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1254__delay_1253__delay_1252__delay_1251___cond_964 <= __delay_data_1253__delay_1252__delay_1251__delay_1250___cond_964;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1271__delay_1270__delay_1269___plus_1025 <= __delay_data_1270__delay_1269__delay_1268___plus_1025;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1289__delay_1288__delay_1287__delay_1286___eq_1031 <= __delay_data_1288__delay_1287__delay_1286__delay_1285___eq_1031;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1318__delay_1317__delay_1316__delay_1315___eq_1034 <= __delay_data_1317__delay_1316__delay_1315__delay_1314___eq_1034;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1238__delay_1237__delay_1236__delay_1235___cond_957 <= __delay_data_1237__delay_1236__delay_1235__delay_1234___cond_957;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1255__delay_1254__delay_1253__delay_1252___cond_964 <= __delay_data_1254__delay_1253__delay_1252__delay_1251___cond_964;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1272__delay_1271__delay_1270___plus_1025 <= __delay_data_1271__delay_1270__delay_1269___plus_1025;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1290__delay_1289__delay_1288__delay_1287___eq_1031 <= __delay_data_1289__delay_1288__delay_1287__delay_1286___eq_1031;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1319__delay_1318__delay_1317__delay_1316___eq_1034 <= __delay_data_1318__delay_1317__delay_1316__delay_1315___eq_1034;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1239__delay_1238__delay_1237__delay_1236___cond_957 <= __delay_data_1238__delay_1237__delay_1236__delay_1235___cond_957;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1256__delay_1255__delay_1254__delay_1253___cond_964 <= __delay_data_1255__delay_1254__delay_1253__delay_1252___cond_964;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1273__delay_1272__delay_1271___plus_1025 <= __delay_data_1272__delay_1271__delay_1270___plus_1025;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1291__delay_1290__delay_1289__delay_1288___eq_1031 <= __delay_data_1290__delay_1289__delay_1288__delay_1287___eq_1031;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1320__delay_1319__delay_1318__delay_1317___eq_1034 <= __delay_data_1319__delay_1318__delay_1317__delay_1316___eq_1034;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1240__delay_1239__delay_1238__delay_1237___cond_957 <= __delay_data_1239__delay_1238__delay_1237__delay_1236___cond_957;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1257__delay_1256__delay_1255__delay_1254___cond_964 <= __delay_data_1256__delay_1255__delay_1254__delay_1253___cond_964;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1274__delay_1273__delay_1272___plus_1025 <= __delay_data_1273__delay_1272__delay_1271___plus_1025;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1292__delay_1291__delay_1290__delay_1289___eq_1031 <= __delay_data_1291__delay_1290__delay_1289__delay_1288___eq_1031;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1321__delay_1320__delay_1319__delay_1318___eq_1034 <= __delay_data_1320__delay_1319__delay_1318__delay_1317___eq_1034;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1241__delay_1240__delay_1239__delay_1238___cond_957 <= __delay_data_1240__delay_1239__delay_1238__delay_1237___cond_957;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1258__delay_1257__delay_1256__delay_1255___cond_964 <= __delay_data_1257__delay_1256__delay_1255__delay_1254___cond_964;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1275__delay_1274__delay_1273___plus_1025 <= __delay_data_1274__delay_1273__delay_1272___plus_1025;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1293__delay_1292__delay_1291__delay_1290___eq_1031 <= __delay_data_1292__delay_1291__delay_1290__delay_1289___eq_1031;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1322__delay_1321__delay_1320__delay_1319___eq_1034 <= __delay_data_1321__delay_1320__delay_1319__delay_1318___eq_1034;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1242__delay_1241__delay_1240__delay_1239___cond_957 <= __delay_data_1241__delay_1240__delay_1239__delay_1238___cond_957;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1259__delay_1258__delay_1257__delay_1256___cond_964 <= __delay_data_1258__delay_1257__delay_1256__delay_1255___cond_964;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1276__delay_1275__delay_1274___plus_1025 <= __delay_data_1275__delay_1274__delay_1273___plus_1025;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1294__delay_1293__delay_1292__delay_1291___eq_1031 <= __delay_data_1293__delay_1292__delay_1291__delay_1290___eq_1031;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1323__delay_1322__delay_1321__delay_1320___eq_1034 <= __delay_data_1322__delay_1321__delay_1320__delay_1319___eq_1034;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1243__delay_1242__delay_1241__delay_1240___cond_957 <= __delay_data_1242__delay_1241__delay_1240__delay_1239___cond_957;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1260__delay_1259__delay_1258__delay_1257___cond_964 <= __delay_data_1259__delay_1258__delay_1257__delay_1256___cond_964;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1277__delay_1276__delay_1275___plus_1025 <= __delay_data_1276__delay_1275__delay_1274___plus_1025;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1295__delay_1294__delay_1293__delay_1292___eq_1031 <= __delay_data_1294__delay_1293__delay_1292__delay_1291___eq_1031;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1324__delay_1323__delay_1322__delay_1321___eq_1034 <= __delay_data_1323__delay_1322__delay_1321__delay_1320___eq_1034;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _plus_data_1023 <= __substreamoutput_data_1021 + __delay_data_1243__delay_1242__delay_1241__delay_1240___cond_957;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1261__delay_1260__delay_1259__delay_1258___cond_964 <= __delay_data_1260__delay_1259__delay_1258__delay_1257___cond_964;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1278__delay_1277__delay_1276___plus_1025 <= __delay_data_1277__delay_1276__delay_1275___plus_1025;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1296__delay_1295__delay_1294__delay_1293___eq_1031 <= __delay_data_1295__delay_1294__delay_1293__delay_1292___eq_1031;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1325__delay_1324__delay_1323__delay_1322___eq_1034 <= __delay_data_1324__delay_1323__delay_1322__delay_1321___eq_1034;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1337__substreamoutput_1022 <= __substreamoutput_data_1022;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1297__delay_1296__delay_1295__delay_1294___eq_1031 <= __delay_data_1296__delay_1295__delay_1294__delay_1293___eq_1031;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1326__delay_1325__delay_1324__delay_1323___eq_1034 <= __delay_data_1325__delay_1324__delay_1323__delay_1322___eq_1034;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1338__delay_1337__substreamoutput_1022 <= __delay_data_1337__substreamoutput_1022;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1298__delay_1297__delay_1296__delay_1295___eq_1031 <= __delay_data_1297__delay_1296__delay_1295__delay_1294___eq_1031;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1327__delay_1326__delay_1325__delay_1324___eq_1034 <= __delay_data_1326__delay_1325__delay_1324__delay_1323___eq_1034;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1339__delay_1338____substreamoutput_1022 <= __delay_data_1338__delay_1337__substreamoutput_1022;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1299__delay_1298__delay_1297__delay_1296___eq_1031 <= __delay_data_1298__delay_1297__delay_1296__delay_1295___eq_1031;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1328__delay_1327__delay_1326__delay_1325___eq_1034 <= __delay_data_1327__delay_1326__delay_1325__delay_1324___eq_1034;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1340__delay_1339____substreamoutput_1022 <= __delay_data_1339__delay_1338____substreamoutput_1022;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1300__delay_1299__delay_1298__delay_1297___eq_1031 <= __delay_data_1299__delay_1298__delay_1297__delay_1296___eq_1031;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1329__delay_1328__delay_1327__delay_1326___eq_1034 <= __delay_data_1328__delay_1327__delay_1326__delay_1325___eq_1034;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1341__delay_1340____substreamoutput_1022 <= __delay_data_1340__delay_1339____substreamoutput_1022;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1301__delay_1300__delay_1299__delay_1298___eq_1031 <= __delay_data_1300__delay_1299__delay_1298__delay_1297___eq_1031;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1330__delay_1329__delay_1328__delay_1327___eq_1034 <= __delay_data_1329__delay_1328__delay_1327__delay_1326___eq_1034;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1342__delay_1341____substreamoutput_1022 <= __delay_data_1341__delay_1340____substreamoutput_1022;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1302__delay_1301__delay_1300__delay_1299___eq_1031 <= __delay_data_1301__delay_1300__delay_1299__delay_1298___eq_1031;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1331__delay_1330__delay_1329__delay_1328___eq_1034 <= __delay_data_1330__delay_1329__delay_1328__delay_1327___eq_1034;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1343__delay_1342____substreamoutput_1022 <= __delay_data_1342__delay_1341____substreamoutput_1022;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1303__delay_1302__delay_1301__delay_1300___eq_1031 <= __delay_data_1302__delay_1301__delay_1300__delay_1299___eq_1031;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1332__delay_1331__delay_1330__delay_1329___eq_1034 <= __delay_data_1331__delay_1330__delay_1329__delay_1328___eq_1034;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1344__delay_1343____substreamoutput_1022 <= __delay_data_1343__delay_1342____substreamoutput_1022;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1304__delay_1303__delay_1302__delay_1301___eq_1031 <= __delay_data_1303__delay_1302__delay_1301__delay_1300___eq_1031;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1333__delay_1332__delay_1331__delay_1330___eq_1034 <= __delay_data_1332__delay_1331__delay_1330__delay_1329___eq_1034;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1345__delay_1344____substreamoutput_1022 <= __delay_data_1344__delay_1343____substreamoutput_1022;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1305__delay_1304__delay_1303__delay_1302___eq_1031 <= __delay_data_1304__delay_1303__delay_1302__delay_1301___eq_1031;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1334__delay_1333__delay_1332__delay_1331___eq_1034 <= __delay_data_1333__delay_1332__delay_1331__delay_1330___eq_1034;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1346__delay_1345____substreamoutput_1022 <= __delay_data_1345__delay_1344____substreamoutput_1022;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _greaterthan_data_1028 <= __substreamoutput_data_1026 > 1'sd0;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1279__substreamoutput_1026 <= __substreamoutput_data_1026;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1306__delay_1305__delay_1304__delay_1303___eq_1031 <= __delay_data_1305__delay_1304__delay_1303__delay_1302___eq_1031;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1335__delay_1334__delay_1333__delay_1332___eq_1034 <= __delay_data_1334__delay_1333__delay_1332__delay_1331___eq_1034;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1347__delay_1346____substreamoutput_1022 <= __delay_data_1346__delay_1345____substreamoutput_1022;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _cond_data_1030 <= (_greaterthan_data_1028)? __delay_data_1279__substreamoutput_1026 : 1'sd0;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1307__delay_1306__delay_1305__delay_1304___eq_1031 <= __delay_data_1306__delay_1305__delay_1304__delay_1303___eq_1031;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1308__delay_1279__substreamoutput_1026 <= __delay_data_1279__substreamoutput_1026;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1336__delay_1335__delay_1334__delay_1333___eq_1034 <= __delay_data_1335__delay_1334__delay_1333__delay_1332___eq_1034;
      end 
      if(_stream_matmul_55_stream_oready) begin
        __delay_data_1348__delay_1347____substreamoutput_1022 <= __delay_data_1347__delay_1346____substreamoutput_1022;
      end 
      if(_set_flag_1656) begin
        _stream_matmul_55_parameter_0_next_parameter_data <= cparam_matmul_55_stream_reduce_size;
      end 
      if(_stream_matmul_55_source_start) begin
        __variable_wdata_936 <= _stream_matmul_55_parameter_0_next_parameter_data;
      end 
      if(_set_flag_1657) begin
        _stream_matmul_55_parameter_1_next_parameter_data <= matmul_55_col_select;
      end 
      if(_stream_matmul_55_source_start) begin
        __variable_wdata_937 <= _stream_matmul_55_parameter_1_next_parameter_data;
      end 
      if(_set_flag_1658) begin
        _stream_matmul_55_parameter_2_next_parameter_data <= matmul_55_row_select_buf;
      end 
      if(_stream_matmul_55_source_start) begin
        __variable_wdata_938 <= _stream_matmul_55_parameter_2_next_parameter_data;
      end 
      if(_set_flag_1659) begin
        _stream_matmul_55_parameter_3_next_parameter_data <= matmul_55_stream_pad_masks;
      end 
      if(_stream_matmul_55_source_start) begin
        __variable_wdata_939 <= _stream_matmul_55_parameter_3_next_parameter_data;
      end 
      if(_set_flag_1660) begin
        _stream_matmul_55_parameter_4_next_parameter_data <= cparam_matmul_55_stream_omit_mask;
      end 
      if(_stream_matmul_55_source_start) begin
        __variable_wdata_940 <= _stream_matmul_55_parameter_4_next_parameter_data;
      end 
      if(_set_flag_1661) begin
        _stream_matmul_55_parameter_6_next_parameter_data <= cparam_matmul_55_bias_scala;
      end 
      if(_stream_matmul_55_source_start) begin
        __variable_wdata_951 <= _stream_matmul_55_parameter_6_next_parameter_data;
      end 
      if(_set_flag_1662) begin
        _stream_matmul_55_source_7_source_mode <= 5'b10;
        _stream_matmul_55_source_7_source_offset <= (cparam_matmul_55_bias_num == 1)? 0 : matmul_55_och_count_buf;
      end 
      if(_set_flag_1662) begin
        _source_stream_matmul_55_source_7_pat_size_0 <= cparam_matmul_55_stream_reduce_size;
        _source_stream_matmul_55_source_7_pat_stride_0 <= 0;
      end 
      if(_set_flag_1662) begin
        _source_stream_matmul_55_source_7_pat_size_1 <= matmul_55_next_stream_num_ops;
        _source_stream_matmul_55_source_7_pat_stride_1 <= (cparam_matmul_55_bias_num == 1)? 0 : 1;
      end 
      if(_set_flag_1662) begin
        _source_stream_matmul_55_source_7_pat_size_2 <= 1;
        _source_stream_matmul_55_source_7_pat_stride_2 <= 0;
      end 
      if(_set_flag_1662) begin
        _source_stream_matmul_55_source_7_pat_size_3 <= 1;
        _source_stream_matmul_55_source_7_pat_stride_3 <= 0;
      end 
      if(_set_flag_1662) begin
        _stream_matmul_55_source_7_source_sel <= 1;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_7_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _stream_matmul_55_source_7_source_offset_buf <= _stream_matmul_55_source_7_source_offset;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_7_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_7_pat_cur_offset_0 <= 0;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_7_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_7_pat_cur_offset_1 <= 0;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_7_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_7_pat_cur_offset_2 <= 0;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_7_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_7_pat_cur_offset_3 <= 0;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_7_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_7_pat_count_0 <= _source_stream_matmul_55_source_7_pat_size_0 - 1;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_7_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_7_pat_count_1 <= _source_stream_matmul_55_source_7_pat_size_1 - 1;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_7_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_7_pat_count_2 <= _source_stream_matmul_55_source_7_pat_size_2 - 1;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_7_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_7_pat_count_3 <= _source_stream_matmul_55_source_7_pat_size_3 - 1;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_7_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_7_pat_size_buf_0 <= _source_stream_matmul_55_source_7_pat_size_0;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_7_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_7_pat_size_buf_1 <= _source_stream_matmul_55_source_7_pat_size_1;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_7_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_7_pat_size_buf_2 <= _source_stream_matmul_55_source_7_pat_size_2;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_7_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_7_pat_size_buf_3 <= _source_stream_matmul_55_source_7_pat_size_3;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_7_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_7_pat_stride_buf_0 <= _source_stream_matmul_55_source_7_pat_stride_0;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_7_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_7_pat_stride_buf_1 <= _source_stream_matmul_55_source_7_pat_stride_1;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_7_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_7_pat_stride_buf_2 <= _source_stream_matmul_55_source_7_pat_stride_2;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_7_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_7_pat_stride_buf_3 <= _source_stream_matmul_55_source_7_pat_stride_3;
      end 
      if(_stream_matmul_55_stream_oready && _stream_matmul_55_source_busy && _stream_matmul_55_is_root) begin
        __variable_wdata_952 <= _stream_matmul_55_source_7_source_ram_rdata;
      end 
      if((_stream_matmul_55_source_7_source_pat_fsm_0 == 1) && _stream_matmul_55_stream_oready) begin
        _stream_matmul_55_source_7_idle <= 0;
        _stream_matmul_55_source_7_source_ram_raddr <= _stream_matmul_55_source_7_source_pat_all_offset;
        _stream_matmul_55_source_7_source_ram_renable <= 1;
      end 
      if((_stream_matmul_55_source_7_source_pat_fsm_0 == 1) && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_7_pat_cur_offset_0 <= _source_stream_matmul_55_source_7_pat_cur_offset_0 + _source_stream_matmul_55_source_7_pat_stride_buf_0;
        _source_stream_matmul_55_source_7_pat_count_0 <= _source_stream_matmul_55_source_7_pat_count_0 - 1;
      end 
      if((_stream_matmul_55_source_7_source_pat_fsm_0 == 1) && (_source_stream_matmul_55_source_7_pat_count_0 == 0) && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_7_pat_cur_offset_0 <= 0;
        _source_stream_matmul_55_source_7_pat_count_0 <= _source_stream_matmul_55_source_7_pat_size_buf_0 - 1;
      end 
      if((_stream_matmul_55_source_7_source_pat_fsm_0 == 1) && (_source_stream_matmul_55_source_7_pat_count_0 == 0) && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_7_pat_cur_offset_1 <= _source_stream_matmul_55_source_7_pat_cur_offset_1 + _source_stream_matmul_55_source_7_pat_stride_buf_1;
        _source_stream_matmul_55_source_7_pat_count_1 <= _source_stream_matmul_55_source_7_pat_count_1 - 1;
      end 
      if((_stream_matmul_55_source_7_source_pat_fsm_0 == 1) && (_source_stream_matmul_55_source_7_pat_count_0 == 0) && (_source_stream_matmul_55_source_7_pat_count_1 == 0) && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_7_pat_cur_offset_1 <= 0;
        _source_stream_matmul_55_source_7_pat_count_1 <= _source_stream_matmul_55_source_7_pat_size_buf_1 - 1;
      end 
      if((_stream_matmul_55_source_7_source_pat_fsm_0 == 1) && ((_source_stream_matmul_55_source_7_pat_count_0 == 0) && (_source_stream_matmul_55_source_7_pat_count_1 == 0)) && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_7_pat_cur_offset_2 <= _source_stream_matmul_55_source_7_pat_cur_offset_2 + _source_stream_matmul_55_source_7_pat_stride_buf_2;
        _source_stream_matmul_55_source_7_pat_count_2 <= _source_stream_matmul_55_source_7_pat_count_2 - 1;
      end 
      if((_stream_matmul_55_source_7_source_pat_fsm_0 == 1) && ((_source_stream_matmul_55_source_7_pat_count_0 == 0) && (_source_stream_matmul_55_source_7_pat_count_1 == 0)) && (_source_stream_matmul_55_source_7_pat_count_2 == 0) && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_7_pat_cur_offset_2 <= 0;
        _source_stream_matmul_55_source_7_pat_count_2 <= _source_stream_matmul_55_source_7_pat_size_buf_2 - 1;
      end 
      if((_stream_matmul_55_source_7_source_pat_fsm_0 == 1) && ((_source_stream_matmul_55_source_7_pat_count_0 == 0) && (_source_stream_matmul_55_source_7_pat_count_1 == 0) && (_source_stream_matmul_55_source_7_pat_count_2 == 0)) && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_7_pat_cur_offset_3 <= _source_stream_matmul_55_source_7_pat_cur_offset_3 + _source_stream_matmul_55_source_7_pat_stride_buf_3;
        _source_stream_matmul_55_source_7_pat_count_3 <= _source_stream_matmul_55_source_7_pat_count_3 - 1;
      end 
      if((_stream_matmul_55_source_7_source_pat_fsm_0 == 1) && ((_source_stream_matmul_55_source_7_pat_count_0 == 0) && (_source_stream_matmul_55_source_7_pat_count_1 == 0) && (_source_stream_matmul_55_source_7_pat_count_2 == 0)) && (_source_stream_matmul_55_source_7_pat_count_3 == 0) && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_7_pat_cur_offset_3 <= 0;
        _source_stream_matmul_55_source_7_pat_count_3 <= _source_stream_matmul_55_source_7_pat_size_buf_3 - 1;
      end 
      if((_stream_matmul_55_source_7_source_pat_fsm_0 == 1) && _stream_matmul_55_source_stop && _stream_matmul_55_stream_oready) begin
        _stream_matmul_55_source_7_source_ram_renable <= 0;
        _stream_matmul_55_source_7_idle <= 1;
      end 
      if((_stream_matmul_55_source_7_source_pat_fsm_0 == 2) && _stream_matmul_55_stream_oready) begin
        _stream_matmul_55_source_7_source_ram_renable <= 0;
        _stream_matmul_55_source_7_idle <= 1;
      end 
      if(_set_flag_1665) begin
        _stream_matmul_55_parameter_8_next_parameter_data <= cparam_matmul_55_scale_scala;
      end 
      if(_stream_matmul_55_source_start) begin
        __variable_wdata_958 <= _stream_matmul_55_parameter_8_next_parameter_data;
      end 
      if(_set_flag_1666) begin
        _stream_matmul_55_source_9_source_mode <= 5'b10;
        _stream_matmul_55_source_9_source_offset <= (cparam_matmul_55_scale_num == 1)? 0 : matmul_55_och_count_buf;
      end 
      if(_set_flag_1666) begin
        _source_stream_matmul_55_source_9_pat_size_0 <= cparam_matmul_55_stream_reduce_size;
        _source_stream_matmul_55_source_9_pat_stride_0 <= 0;
      end 
      if(_set_flag_1666) begin
        _source_stream_matmul_55_source_9_pat_size_1 <= matmul_55_next_stream_num_ops;
        _source_stream_matmul_55_source_9_pat_stride_1 <= (cparam_matmul_55_scale_num == 1)? 0 : 1;
      end 
      if(_set_flag_1666) begin
        _source_stream_matmul_55_source_9_pat_size_2 <= 1;
        _source_stream_matmul_55_source_9_pat_stride_2 <= 0;
      end 
      if(_set_flag_1666) begin
        _source_stream_matmul_55_source_9_pat_size_3 <= 1;
        _source_stream_matmul_55_source_9_pat_stride_3 <= 0;
      end 
      if(_set_flag_1666) begin
        _stream_matmul_55_source_9_source_sel <= 2;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_9_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _stream_matmul_55_source_9_source_offset_buf <= _stream_matmul_55_source_9_source_offset;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_9_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_9_pat_cur_offset_0 <= 0;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_9_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_9_pat_cur_offset_1 <= 0;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_9_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_9_pat_cur_offset_2 <= 0;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_9_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_9_pat_cur_offset_3 <= 0;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_9_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_9_pat_count_0 <= _source_stream_matmul_55_source_9_pat_size_0 - 1;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_9_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_9_pat_count_1 <= _source_stream_matmul_55_source_9_pat_size_1 - 1;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_9_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_9_pat_count_2 <= _source_stream_matmul_55_source_9_pat_size_2 - 1;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_9_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_9_pat_count_3 <= _source_stream_matmul_55_source_9_pat_size_3 - 1;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_9_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_9_pat_size_buf_0 <= _source_stream_matmul_55_source_9_pat_size_0;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_9_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_9_pat_size_buf_1 <= _source_stream_matmul_55_source_9_pat_size_1;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_9_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_9_pat_size_buf_2 <= _source_stream_matmul_55_source_9_pat_size_2;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_9_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_9_pat_size_buf_3 <= _source_stream_matmul_55_source_9_pat_size_3;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_9_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_9_pat_stride_buf_0 <= _source_stream_matmul_55_source_9_pat_stride_0;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_9_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_9_pat_stride_buf_1 <= _source_stream_matmul_55_source_9_pat_stride_1;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_9_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_9_pat_stride_buf_2 <= _source_stream_matmul_55_source_9_pat_stride_2;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_9_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_9_pat_stride_buf_3 <= _source_stream_matmul_55_source_9_pat_stride_3;
      end 
      if(_stream_matmul_55_stream_oready && _stream_matmul_55_source_busy && _stream_matmul_55_is_root) begin
        __variable_wdata_959 <= _stream_matmul_55_source_9_source_ram_rdata;
      end 
      if((_stream_matmul_55_source_9_source_pat_fsm_1 == 1) && _stream_matmul_55_stream_oready) begin
        _stream_matmul_55_source_9_idle <= 0;
        _stream_matmul_55_source_9_source_ram_raddr <= _stream_matmul_55_source_9_source_pat_all_offset;
        _stream_matmul_55_source_9_source_ram_renable <= 1;
      end 
      if((_stream_matmul_55_source_9_source_pat_fsm_1 == 1) && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_9_pat_cur_offset_0 <= _source_stream_matmul_55_source_9_pat_cur_offset_0 + _source_stream_matmul_55_source_9_pat_stride_buf_0;
        _source_stream_matmul_55_source_9_pat_count_0 <= _source_stream_matmul_55_source_9_pat_count_0 - 1;
      end 
      if((_stream_matmul_55_source_9_source_pat_fsm_1 == 1) && (_source_stream_matmul_55_source_9_pat_count_0 == 0) && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_9_pat_cur_offset_0 <= 0;
        _source_stream_matmul_55_source_9_pat_count_0 <= _source_stream_matmul_55_source_9_pat_size_buf_0 - 1;
      end 
      if((_stream_matmul_55_source_9_source_pat_fsm_1 == 1) && (_source_stream_matmul_55_source_9_pat_count_0 == 0) && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_9_pat_cur_offset_1 <= _source_stream_matmul_55_source_9_pat_cur_offset_1 + _source_stream_matmul_55_source_9_pat_stride_buf_1;
        _source_stream_matmul_55_source_9_pat_count_1 <= _source_stream_matmul_55_source_9_pat_count_1 - 1;
      end 
      if((_stream_matmul_55_source_9_source_pat_fsm_1 == 1) && (_source_stream_matmul_55_source_9_pat_count_0 == 0) && (_source_stream_matmul_55_source_9_pat_count_1 == 0) && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_9_pat_cur_offset_1 <= 0;
        _source_stream_matmul_55_source_9_pat_count_1 <= _source_stream_matmul_55_source_9_pat_size_buf_1 - 1;
      end 
      if((_stream_matmul_55_source_9_source_pat_fsm_1 == 1) && ((_source_stream_matmul_55_source_9_pat_count_0 == 0) && (_source_stream_matmul_55_source_9_pat_count_1 == 0)) && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_9_pat_cur_offset_2 <= _source_stream_matmul_55_source_9_pat_cur_offset_2 + _source_stream_matmul_55_source_9_pat_stride_buf_2;
        _source_stream_matmul_55_source_9_pat_count_2 <= _source_stream_matmul_55_source_9_pat_count_2 - 1;
      end 
      if((_stream_matmul_55_source_9_source_pat_fsm_1 == 1) && ((_source_stream_matmul_55_source_9_pat_count_0 == 0) && (_source_stream_matmul_55_source_9_pat_count_1 == 0)) && (_source_stream_matmul_55_source_9_pat_count_2 == 0) && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_9_pat_cur_offset_2 <= 0;
        _source_stream_matmul_55_source_9_pat_count_2 <= _source_stream_matmul_55_source_9_pat_size_buf_2 - 1;
      end 
      if((_stream_matmul_55_source_9_source_pat_fsm_1 == 1) && ((_source_stream_matmul_55_source_9_pat_count_0 == 0) && (_source_stream_matmul_55_source_9_pat_count_1 == 0) && (_source_stream_matmul_55_source_9_pat_count_2 == 0)) && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_9_pat_cur_offset_3 <= _source_stream_matmul_55_source_9_pat_cur_offset_3 + _source_stream_matmul_55_source_9_pat_stride_buf_3;
        _source_stream_matmul_55_source_9_pat_count_3 <= _source_stream_matmul_55_source_9_pat_count_3 - 1;
      end 
      if((_stream_matmul_55_source_9_source_pat_fsm_1 == 1) && ((_source_stream_matmul_55_source_9_pat_count_0 == 0) && (_source_stream_matmul_55_source_9_pat_count_1 == 0) && (_source_stream_matmul_55_source_9_pat_count_2 == 0)) && (_source_stream_matmul_55_source_9_pat_count_3 == 0) && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_9_pat_cur_offset_3 <= 0;
        _source_stream_matmul_55_source_9_pat_count_3 <= _source_stream_matmul_55_source_9_pat_size_buf_3 - 1;
      end 
      if((_stream_matmul_55_source_9_source_pat_fsm_1 == 1) && _stream_matmul_55_source_stop && _stream_matmul_55_stream_oready) begin
        _stream_matmul_55_source_9_source_ram_renable <= 0;
        _stream_matmul_55_source_9_idle <= 1;
      end 
      if((_stream_matmul_55_source_9_source_pat_fsm_1 == 2) && _stream_matmul_55_stream_oready) begin
        _stream_matmul_55_source_9_source_ram_renable <= 0;
        _stream_matmul_55_source_9_idle <= 1;
      end 
      if(_set_flag_1679) begin
        _stream_matmul_55_parameter_10_next_parameter_data <= 1;
      end 
      if(_stream_matmul_55_source_start) begin
        __variable_wdata_965 <= _stream_matmul_55_parameter_10_next_parameter_data;
      end 
      if(_set_flag_1680) begin
        _stream_matmul_55_source_11_source_mode <= 5'b0;
        _stream_matmul_55_source_11_source_empty_data <= 0;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_stream_oready && !(|(_stream_matmul_55_source_11_source_mode & 5'b0))) begin
        _stream_matmul_55_source_11_idle <= 1;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_stream_oready && !(|(_stream_matmul_55_source_11_source_mode & 5'b0)) && _stream_matmul_55_is_root) begin
        __variable_wdata_966 <= _stream_matmul_55_source_11_source_empty_data;
      end 
      if(_set_flag_1681) begin
        _stream_matmul_55_parameter_12_next_parameter_data <= 1;
      end 
      if(_stream_matmul_55_source_start) begin
        __variable_wdata_972 <= _stream_matmul_55_parameter_12_next_parameter_data;
      end 
      if(_set_flag_1682) begin
        _stream_matmul_55_source_13_source_mode <= 5'b0;
        _stream_matmul_55_source_13_source_empty_data <= 0;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_stream_oready && !(|(_stream_matmul_55_source_13_source_mode & 5'b0))) begin
        _stream_matmul_55_source_13_idle <= 1;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_stream_oready && !(|(_stream_matmul_55_source_13_source_mode & 5'b0)) && _stream_matmul_55_is_root) begin
        __variable_wdata_973 <= _stream_matmul_55_source_13_source_empty_data;
      end 
      if(_set_flag_1683) begin
        _stream_matmul_55_parameter_14_next_parameter_data <= 1;
      end 
      if(_stream_matmul_55_source_start) begin
        __variable_wdata_979 <= _stream_matmul_55_parameter_14_next_parameter_data;
      end 
      if(_set_flag_1684) begin
        _stream_matmul_55_source_15_source_mode <= 5'b0;
        _stream_matmul_55_source_15_source_empty_data <= 0;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_stream_oready && !(|(_stream_matmul_55_source_15_source_mode & 5'b0))) begin
        _stream_matmul_55_source_15_idle <= 1;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_stream_oready && !(|(_stream_matmul_55_source_15_source_mode & 5'b0)) && _stream_matmul_55_is_root) begin
        __variable_wdata_980 <= _stream_matmul_55_source_15_source_empty_data;
      end 
      if(_set_flag_1685) begin
        _stream_matmul_55_parameter_16_next_parameter_data <= cparam_matmul_55_cshamt_mul_value;
      end 
      if(_stream_matmul_55_source_start) begin
        __variable_wdata_986 <= _stream_matmul_55_parameter_16_next_parameter_data;
      end 
      if(_set_flag_1686) begin
        _stream_matmul_55_parameter_17_next_parameter_data <= cparam_matmul_55_cshamt_sum_value;
      end 
      if(_stream_matmul_55_source_start) begin
        __variable_wdata_987 <= _stream_matmul_55_parameter_17_next_parameter_data;
      end 
      if(_set_flag_1687) begin
        _stream_matmul_55_parameter_18_next_parameter_data <= cparam_matmul_55_cshamt_out_value;
      end 
      if(_stream_matmul_55_source_start) begin
        __variable_wdata_988 <= _stream_matmul_55_parameter_18_next_parameter_data;
      end 
      if(_set_flag_1688) begin
        _stream_matmul_55_parameter_19_next_parameter_data <= cparam_matmul_55_act_func_index;
      end 
      if(_stream_matmul_55_source_start) begin
        __variable_wdata_989 <= _stream_matmul_55_parameter_19_next_parameter_data;
      end 
      if(_set_flag_1689) begin
        _stream_matmul_55_source_20_source_mode <= 5'b10;
        _stream_matmul_55_source_20_source_offset <= matmul_55_stream_act_local_0 + matmul_55_act_page_comp_offset_buf_0;
      end 
      if(_set_flag_1689) begin
        _source_stream_matmul_55_source_20_pat_size_0 <= cparam_matmul_55_stream_reduce_size;
        _source_stream_matmul_55_source_20_pat_stride_0 <= 1;
      end 
      if(_set_flag_1689) begin
        _source_stream_matmul_55_source_20_pat_size_1 <= matmul_55_next_stream_num_ops;
        _source_stream_matmul_55_source_20_pat_stride_1 <= 0;
      end 
      if(_set_flag_1689) begin
        _source_stream_matmul_55_source_20_pat_size_2 <= 1;
        _source_stream_matmul_55_source_20_pat_stride_2 <= 0;
      end 
      if(_set_flag_1689) begin
        _source_stream_matmul_55_source_20_pat_size_3 <= 1;
        _source_stream_matmul_55_source_20_pat_stride_3 <= 0;
      end 
      if(_set_flag_1689) begin
        _stream_matmul_55_source_20_source_sel <= 3;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_20_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _stream_matmul_55_source_20_source_offset_buf <= _stream_matmul_55_source_20_source_offset;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_20_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_20_pat_cur_offset_0 <= 0;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_20_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_20_pat_cur_offset_1 <= 0;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_20_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_20_pat_cur_offset_2 <= 0;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_20_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_20_pat_cur_offset_3 <= 0;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_20_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_20_pat_count_0 <= _source_stream_matmul_55_source_20_pat_size_0 - 1;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_20_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_20_pat_count_1 <= _source_stream_matmul_55_source_20_pat_size_1 - 1;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_20_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_20_pat_count_2 <= _source_stream_matmul_55_source_20_pat_size_2 - 1;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_20_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_20_pat_count_3 <= _source_stream_matmul_55_source_20_pat_size_3 - 1;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_20_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_20_pat_size_buf_0 <= _source_stream_matmul_55_source_20_pat_size_0;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_20_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_20_pat_size_buf_1 <= _source_stream_matmul_55_source_20_pat_size_1;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_20_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_20_pat_size_buf_2 <= _source_stream_matmul_55_source_20_pat_size_2;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_20_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_20_pat_size_buf_3 <= _source_stream_matmul_55_source_20_pat_size_3;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_20_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_20_pat_stride_buf_0 <= _source_stream_matmul_55_source_20_pat_stride_0;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_20_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_20_pat_stride_buf_1 <= _source_stream_matmul_55_source_20_pat_stride_1;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_20_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_20_pat_stride_buf_2 <= _source_stream_matmul_55_source_20_pat_stride_2;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_20_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_20_pat_stride_buf_3 <= _source_stream_matmul_55_source_20_pat_stride_3;
      end 
      if(_stream_matmul_55_stream_oready && _stream_matmul_55_source_busy && _stream_matmul_55_is_root) begin
        __variable_wdata_990 <= _stream_matmul_55_source_20_source_ram_rdata;
      end 
      if((_stream_matmul_55_source_20_source_pat_fsm_2 == 1) && _stream_matmul_55_stream_oready) begin
        _stream_matmul_55_source_20_idle <= 0;
        _stream_matmul_55_source_20_source_ram_raddr <= _stream_matmul_55_source_20_source_pat_all_offset;
        _stream_matmul_55_source_20_source_ram_renable <= 1;
      end 
      if((_stream_matmul_55_source_20_source_pat_fsm_2 == 1) && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_20_pat_cur_offset_0 <= _source_stream_matmul_55_source_20_pat_cur_offset_0 + _source_stream_matmul_55_source_20_pat_stride_buf_0;
        _source_stream_matmul_55_source_20_pat_count_0 <= _source_stream_matmul_55_source_20_pat_count_0 - 1;
      end 
      if((_stream_matmul_55_source_20_source_pat_fsm_2 == 1) && (_source_stream_matmul_55_source_20_pat_count_0 == 0) && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_20_pat_cur_offset_0 <= 0;
        _source_stream_matmul_55_source_20_pat_count_0 <= _source_stream_matmul_55_source_20_pat_size_buf_0 - 1;
      end 
      if((_stream_matmul_55_source_20_source_pat_fsm_2 == 1) && (_source_stream_matmul_55_source_20_pat_count_0 == 0) && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_20_pat_cur_offset_1 <= _source_stream_matmul_55_source_20_pat_cur_offset_1 + _source_stream_matmul_55_source_20_pat_stride_buf_1;
        _source_stream_matmul_55_source_20_pat_count_1 <= _source_stream_matmul_55_source_20_pat_count_1 - 1;
      end 
      if((_stream_matmul_55_source_20_source_pat_fsm_2 == 1) && (_source_stream_matmul_55_source_20_pat_count_0 == 0) && (_source_stream_matmul_55_source_20_pat_count_1 == 0) && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_20_pat_cur_offset_1 <= 0;
        _source_stream_matmul_55_source_20_pat_count_1 <= _source_stream_matmul_55_source_20_pat_size_buf_1 - 1;
      end 
      if((_stream_matmul_55_source_20_source_pat_fsm_2 == 1) && ((_source_stream_matmul_55_source_20_pat_count_0 == 0) && (_source_stream_matmul_55_source_20_pat_count_1 == 0)) && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_20_pat_cur_offset_2 <= _source_stream_matmul_55_source_20_pat_cur_offset_2 + _source_stream_matmul_55_source_20_pat_stride_buf_2;
        _source_stream_matmul_55_source_20_pat_count_2 <= _source_stream_matmul_55_source_20_pat_count_2 - 1;
      end 
      if((_stream_matmul_55_source_20_source_pat_fsm_2 == 1) && ((_source_stream_matmul_55_source_20_pat_count_0 == 0) && (_source_stream_matmul_55_source_20_pat_count_1 == 0)) && (_source_stream_matmul_55_source_20_pat_count_2 == 0) && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_20_pat_cur_offset_2 <= 0;
        _source_stream_matmul_55_source_20_pat_count_2 <= _source_stream_matmul_55_source_20_pat_size_buf_2 - 1;
      end 
      if((_stream_matmul_55_source_20_source_pat_fsm_2 == 1) && ((_source_stream_matmul_55_source_20_pat_count_0 == 0) && (_source_stream_matmul_55_source_20_pat_count_1 == 0) && (_source_stream_matmul_55_source_20_pat_count_2 == 0)) && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_20_pat_cur_offset_3 <= _source_stream_matmul_55_source_20_pat_cur_offset_3 + _source_stream_matmul_55_source_20_pat_stride_buf_3;
        _source_stream_matmul_55_source_20_pat_count_3 <= _source_stream_matmul_55_source_20_pat_count_3 - 1;
      end 
      if((_stream_matmul_55_source_20_source_pat_fsm_2 == 1) && ((_source_stream_matmul_55_source_20_pat_count_0 == 0) && (_source_stream_matmul_55_source_20_pat_count_1 == 0) && (_source_stream_matmul_55_source_20_pat_count_2 == 0)) && (_source_stream_matmul_55_source_20_pat_count_3 == 0) && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_20_pat_cur_offset_3 <= 0;
        _source_stream_matmul_55_source_20_pat_count_3 <= _source_stream_matmul_55_source_20_pat_size_buf_3 - 1;
      end 
      if((_stream_matmul_55_source_20_source_pat_fsm_2 == 1) && _stream_matmul_55_source_stop && _stream_matmul_55_stream_oready) begin
        _stream_matmul_55_source_20_source_ram_renable <= 0;
        _stream_matmul_55_source_20_idle <= 1;
      end 
      if((_stream_matmul_55_source_20_source_pat_fsm_2 == 2) && _stream_matmul_55_stream_oready) begin
        _stream_matmul_55_source_20_source_ram_renable <= 0;
        _stream_matmul_55_source_20_idle <= 1;
      end 
      if(_set_flag_1702) begin
        _stream_matmul_55_source_21_source_mode <= 5'b10;
        _stream_matmul_55_source_21_source_offset <= matmul_55_filter_page_comp_offset_buf;
      end 
      if(_set_flag_1702) begin
        _source_stream_matmul_55_source_21_pat_size_0 <= cparam_matmul_55_stream_reduce_size;
        _source_stream_matmul_55_source_21_pat_stride_0 <= 1;
      end 
      if(_set_flag_1702) begin
        _source_stream_matmul_55_source_21_pat_size_1 <= matmul_55_next_stream_num_ops;
        _source_stream_matmul_55_source_21_pat_stride_1 <= cparam_matmul_55_stream_aligned_reduce_size;
      end 
      if(_set_flag_1702) begin
        _source_stream_matmul_55_source_21_pat_size_2 <= 1;
        _source_stream_matmul_55_source_21_pat_stride_2 <= 0;
      end 
      if(_set_flag_1702) begin
        _source_stream_matmul_55_source_21_pat_size_3 <= 1;
        _source_stream_matmul_55_source_21_pat_stride_3 <= 0;
      end 
      if(_set_flag_1702) begin
        _stream_matmul_55_source_21_source_sel <= 4;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_21_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _stream_matmul_55_source_21_source_offset_buf <= _stream_matmul_55_source_21_source_offset;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_21_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_21_pat_cur_offset_0 <= 0;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_21_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_21_pat_cur_offset_1 <= 0;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_21_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_21_pat_cur_offset_2 <= 0;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_21_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_21_pat_cur_offset_3 <= 0;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_21_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_21_pat_count_0 <= _source_stream_matmul_55_source_21_pat_size_0 - 1;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_21_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_21_pat_count_1 <= _source_stream_matmul_55_source_21_pat_size_1 - 1;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_21_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_21_pat_count_2 <= _source_stream_matmul_55_source_21_pat_size_2 - 1;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_21_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_21_pat_count_3 <= _source_stream_matmul_55_source_21_pat_size_3 - 1;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_21_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_21_pat_size_buf_0 <= _source_stream_matmul_55_source_21_pat_size_0;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_21_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_21_pat_size_buf_1 <= _source_stream_matmul_55_source_21_pat_size_1;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_21_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_21_pat_size_buf_2 <= _source_stream_matmul_55_source_21_pat_size_2;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_21_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_21_pat_size_buf_3 <= _source_stream_matmul_55_source_21_pat_size_3;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_21_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_21_pat_stride_buf_0 <= _source_stream_matmul_55_source_21_pat_stride_0;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_21_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_21_pat_stride_buf_1 <= _source_stream_matmul_55_source_21_pat_stride_1;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_21_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_21_pat_stride_buf_2 <= _source_stream_matmul_55_source_21_pat_stride_2;
      end 
      if(_stream_matmul_55_source_start && _stream_matmul_55_source_21_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_21_pat_stride_buf_3 <= _source_stream_matmul_55_source_21_pat_stride_3;
      end 
      if(_stream_matmul_55_stream_oready && _stream_matmul_55_source_busy && _stream_matmul_55_is_root) begin
        __variable_wdata_1004 <= _stream_matmul_55_source_21_source_ram_rdata;
      end 
      if((_stream_matmul_55_source_21_source_pat_fsm_3 == 1) && _stream_matmul_55_stream_oready) begin
        _stream_matmul_55_source_21_idle <= 0;
        _stream_matmul_55_source_21_source_ram_raddr <= _stream_matmul_55_source_21_source_pat_all_offset;
        _stream_matmul_55_source_21_source_ram_renable <= 1;
      end 
      if((_stream_matmul_55_source_21_source_pat_fsm_3 == 1) && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_21_pat_cur_offset_0 <= _source_stream_matmul_55_source_21_pat_cur_offset_0 + _source_stream_matmul_55_source_21_pat_stride_buf_0;
        _source_stream_matmul_55_source_21_pat_count_0 <= _source_stream_matmul_55_source_21_pat_count_0 - 1;
      end 
      if((_stream_matmul_55_source_21_source_pat_fsm_3 == 1) && (_source_stream_matmul_55_source_21_pat_count_0 == 0) && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_21_pat_cur_offset_0 <= 0;
        _source_stream_matmul_55_source_21_pat_count_0 <= _source_stream_matmul_55_source_21_pat_size_buf_0 - 1;
      end 
      if((_stream_matmul_55_source_21_source_pat_fsm_3 == 1) && (_source_stream_matmul_55_source_21_pat_count_0 == 0) && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_21_pat_cur_offset_1 <= _source_stream_matmul_55_source_21_pat_cur_offset_1 + _source_stream_matmul_55_source_21_pat_stride_buf_1;
        _source_stream_matmul_55_source_21_pat_count_1 <= _source_stream_matmul_55_source_21_pat_count_1 - 1;
      end 
      if((_stream_matmul_55_source_21_source_pat_fsm_3 == 1) && (_source_stream_matmul_55_source_21_pat_count_0 == 0) && (_source_stream_matmul_55_source_21_pat_count_1 == 0) && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_21_pat_cur_offset_1 <= 0;
        _source_stream_matmul_55_source_21_pat_count_1 <= _source_stream_matmul_55_source_21_pat_size_buf_1 - 1;
      end 
      if((_stream_matmul_55_source_21_source_pat_fsm_3 == 1) && ((_source_stream_matmul_55_source_21_pat_count_0 == 0) && (_source_stream_matmul_55_source_21_pat_count_1 == 0)) && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_21_pat_cur_offset_2 <= _source_stream_matmul_55_source_21_pat_cur_offset_2 + _source_stream_matmul_55_source_21_pat_stride_buf_2;
        _source_stream_matmul_55_source_21_pat_count_2 <= _source_stream_matmul_55_source_21_pat_count_2 - 1;
      end 
      if((_stream_matmul_55_source_21_source_pat_fsm_3 == 1) && ((_source_stream_matmul_55_source_21_pat_count_0 == 0) && (_source_stream_matmul_55_source_21_pat_count_1 == 0)) && (_source_stream_matmul_55_source_21_pat_count_2 == 0) && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_21_pat_cur_offset_2 <= 0;
        _source_stream_matmul_55_source_21_pat_count_2 <= _source_stream_matmul_55_source_21_pat_size_buf_2 - 1;
      end 
      if((_stream_matmul_55_source_21_source_pat_fsm_3 == 1) && ((_source_stream_matmul_55_source_21_pat_count_0 == 0) && (_source_stream_matmul_55_source_21_pat_count_1 == 0) && (_source_stream_matmul_55_source_21_pat_count_2 == 0)) && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_21_pat_cur_offset_3 <= _source_stream_matmul_55_source_21_pat_cur_offset_3 + _source_stream_matmul_55_source_21_pat_stride_buf_3;
        _source_stream_matmul_55_source_21_pat_count_3 <= _source_stream_matmul_55_source_21_pat_count_3 - 1;
      end 
      if((_stream_matmul_55_source_21_source_pat_fsm_3 == 1) && ((_source_stream_matmul_55_source_21_pat_count_0 == 0) && (_source_stream_matmul_55_source_21_pat_count_1 == 0) && (_source_stream_matmul_55_source_21_pat_count_2 == 0)) && (_source_stream_matmul_55_source_21_pat_count_3 == 0) && _stream_matmul_55_stream_oready) begin
        _source_stream_matmul_55_source_21_pat_cur_offset_3 <= 0;
        _source_stream_matmul_55_source_21_pat_count_3 <= _source_stream_matmul_55_source_21_pat_size_buf_3 - 1;
      end 
      if((_stream_matmul_55_source_21_source_pat_fsm_3 == 1) && _stream_matmul_55_source_stop && _stream_matmul_55_stream_oready) begin
        _stream_matmul_55_source_21_source_ram_renable <= 0;
        _stream_matmul_55_source_21_idle <= 1;
      end 
      if((_stream_matmul_55_source_21_source_pat_fsm_3 == 2) && _stream_matmul_55_stream_oready) begin
        _stream_matmul_55_source_21_source_ram_renable <= 0;
        _stream_matmul_55_source_21_idle <= 1;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1716 <= _set_flag_1715;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1717 <= _tmp_1716;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1718 <= _tmp_1717;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1719 <= _tmp_1718;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1720 <= _tmp_1719;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1721 <= _tmp_1720;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1722 <= _tmp_1721;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1723 <= _tmp_1722;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1724 <= _tmp_1723;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1725 <= _tmp_1724;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1726 <= _tmp_1725;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1727 <= _tmp_1726;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1728 <= _tmp_1727;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1729 <= _tmp_1728;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1730 <= _tmp_1729;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1731 <= _tmp_1730;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1732 <= _tmp_1731;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1733 <= _tmp_1732;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1734 <= _tmp_1733;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1735 <= _tmp_1734;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1736 <= _tmp_1735;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1737 <= _tmp_1736;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1738 <= _tmp_1737;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1739 <= _tmp_1738;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1740 <= _tmp_1739;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1741 <= _tmp_1740;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1742 <= _tmp_1741;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1743 <= _tmp_1742;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1744 <= _tmp_1743;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1745 <= _tmp_1744;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1746 <= _tmp_1745;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1749 <= _tmp_1748;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1750 <= _tmp_1749;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1751 <= _tmp_1750;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1752 <= _tmp_1751;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1753 <= _tmp_1752;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1754 <= _tmp_1753;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1755 <= _tmp_1754;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1756 <= _tmp_1755;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1757 <= _tmp_1756;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1758 <= _tmp_1757;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1759 <= _tmp_1758;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1760 <= _tmp_1759;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1761 <= _tmp_1760;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1762 <= _tmp_1761;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1763 <= _tmp_1762;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1764 <= _tmp_1763;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1765 <= _tmp_1764;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1766 <= _tmp_1765;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1767 <= _tmp_1766;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1768 <= _tmp_1767;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1769 <= _tmp_1768;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1770 <= _tmp_1769;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1771 <= _tmp_1770;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1772 <= _tmp_1771;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1773 <= _tmp_1772;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1774 <= _tmp_1773;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1775 <= _tmp_1774;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1776 <= _tmp_1775;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1777 <= _tmp_1776;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1778 <= _tmp_1777;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1779 <= _tmp_1778;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1780 <= matmul_55_next_stream_num_ops;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1781 <= _tmp_1780;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1782 <= _tmp_1781;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1783 <= _tmp_1782;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1784 <= _tmp_1783;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1785 <= _tmp_1784;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1786 <= _tmp_1785;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1787 <= _tmp_1786;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1788 <= _tmp_1787;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1789 <= _tmp_1788;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1790 <= _tmp_1789;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1791 <= _tmp_1790;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1792 <= _tmp_1791;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1793 <= _tmp_1792;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1794 <= _tmp_1793;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1795 <= _tmp_1794;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1796 <= _tmp_1795;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1797 <= _tmp_1796;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1798 <= _tmp_1797;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1799 <= _tmp_1798;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1800 <= _tmp_1799;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1801 <= _tmp_1800;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1802 <= _tmp_1801;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1803 <= _tmp_1802;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1804 <= _tmp_1803;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1805 <= _tmp_1804;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1806 <= _tmp_1805;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1807 <= _tmp_1806;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1808 <= _tmp_1807;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1809 <= _tmp_1808;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1810 <= _tmp_1809;
      end 
      if(_tmp_1746) begin
        _stream_matmul_55_sink_26_sink_mode <= 5'b1;
        _stream_matmul_55_sink_26_sink_offset <= _tmp_1779;
        _stream_matmul_55_sink_26_sink_size <= _tmp_1810;
        _stream_matmul_55_sink_26_sink_stride <= 1;
      end 
      if(_tmp_1746) begin
        _stream_matmul_55_sink_26_sink_sel <= 5;
      end 
      if(_stream_matmul_55_sink_start && _stream_matmul_55_sink_26_sink_mode & 5'b1 && _stream_matmul_55_stream_oready) begin
        _stream_matmul_55_sink_26_sink_offset_buf <= _stream_matmul_55_sink_26_sink_offset;
        _stream_matmul_55_sink_26_sink_size_buf <= _stream_matmul_55_sink_26_sink_size;
        _stream_matmul_55_sink_26_sink_stride_buf <= _stream_matmul_55_sink_26_sink_stride;
      end 
      if((_stream_matmul_55_sink_26_sink_fsm_4 == 1) && _stream_matmul_55_stream_oready) begin
        _stream_matmul_55_sink_26_sink_waddr <= _stream_matmul_55_sink_26_sink_offset_buf - _stream_matmul_55_sink_26_sink_stride_buf;
        _stream_matmul_55_sink_26_sink_count <= _stream_matmul_55_sink_26_sink_size_buf;
      end 
      if((_stream_matmul_55_sink_26_sink_fsm_4 == 2) && stream_matmul_55_sink_27_data && _stream_matmul_55_stream_oready) begin
        _stream_matmul_55_sink_26_sink_waddr <= _stream_matmul_55_sink_26_sink_waddr + _stream_matmul_55_sink_26_sink_stride_buf;
        _stream_matmul_55_sink_26_sink_wdata <= stream_matmul_55_sink_26_data;
        _stream_matmul_55_sink_26_sink_wenable <= 1;
        _stream_matmul_55_sink_26_sink_count <= _stream_matmul_55_sink_26_sink_count - 1;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1823 <= _stream_matmul_55_source_start;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1824 <= _tmp_1823;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1825 <= _tmp_1824;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1826 <= _stream_matmul_55_source_start;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1827 <= _tmp_1826;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1828 <= _tmp_1827;
      end 
      if(_stream_matmul_55_stream_oready && _tmp_1828) begin
        __variable_wdata_941 <= 1;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1829 <= _stream_matmul_55_source_start;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1830 <= _tmp_1829;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1831 <= _tmp_1830;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1832 <= _tmp_1831;
      end 
      if(_stream_matmul_55_stream_oready && _tmp_1832) begin
        __variable_wdata_941 <= 0;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1835 <= _tmp_1834;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1838 <= _tmp_1837;
      end 
      if(_stream_matmul_55_stream_oready && _tmp_1838) begin
        __variable_wdata_941 <= 1;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1839 <= _stream_matmul_55_source_start;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1840 <= _tmp_1839;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1841 <= _tmp_1840;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1842 <= _tmp_1841;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1843 <= _tmp_1842;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1844 <= _tmp_1843;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1845 <= _tmp_1844;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1846 <= _tmp_1845;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1847 <= _tmp_1846;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1848 <= _tmp_1847;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1849 <= _tmp_1848;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1850 <= _tmp_1849;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1851 <= _tmp_1850;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1852 <= _tmp_1851;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1853 <= _tmp_1852;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1854 <= _tmp_1853;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1855 <= _tmp_1854;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1856 <= _tmp_1855;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1857 <= _tmp_1856;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1858 <= _tmp_1857;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1859 <= _tmp_1858;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1860 <= _tmp_1859;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1861 <= _tmp_1860;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1862 <= _tmp_1861;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1863 <= _tmp_1862;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1864 <= _tmp_1863;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1865 <= _tmp_1864;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1866 <= _tmp_1865;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1867 <= _tmp_1866;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1868 <= _tmp_1867;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1869 <= _tmp_1868;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1870 <= _stream_matmul_55_source_stop;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1871 <= _tmp_1870;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1872 <= _tmp_1871;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1873 <= _tmp_1872;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1874 <= _tmp_1873;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1875 <= _tmp_1874;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1876 <= _tmp_1875;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1877 <= _tmp_1876;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1878 <= _tmp_1877;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1879 <= _tmp_1878;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1880 <= _tmp_1879;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1881 <= _tmp_1880;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1882 <= _tmp_1881;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1883 <= _tmp_1882;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1884 <= _tmp_1883;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1885 <= _tmp_1884;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1886 <= _tmp_1885;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1887 <= _tmp_1886;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1888 <= _tmp_1887;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1889 <= _tmp_1888;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1890 <= _tmp_1889;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1891 <= _tmp_1890;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1892 <= _tmp_1891;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1893 <= _tmp_1892;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1894 <= _tmp_1893;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1895 <= _tmp_1894;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1896 <= _tmp_1895;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1897 <= _tmp_1896;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1898 <= _tmp_1897;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1899 <= _tmp_1898;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1900 <= _tmp_1899;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1901 <= _stream_matmul_55_source_busy;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1902 <= _tmp_1901;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1903 <= _tmp_1902;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1904 <= _tmp_1903;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1905 <= _tmp_1904;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1906 <= _tmp_1905;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1907 <= _tmp_1906;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1908 <= _tmp_1907;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1909 <= _tmp_1908;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1910 <= _tmp_1909;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1911 <= _tmp_1910;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1912 <= _tmp_1911;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1913 <= _tmp_1912;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1914 <= _tmp_1913;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1915 <= _tmp_1914;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1916 <= _tmp_1915;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1917 <= _tmp_1916;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1918 <= _tmp_1917;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1919 <= _tmp_1918;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1920 <= _tmp_1919;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1921 <= _tmp_1920;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1922 <= _tmp_1921;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1923 <= _tmp_1922;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1924 <= _tmp_1923;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1925 <= _tmp_1924;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1926 <= _tmp_1925;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1927 <= _tmp_1926;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1928 <= _tmp_1927;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1929 <= _tmp_1928;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1930 <= _tmp_1929;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1931 <= _tmp_1930;
      end 
      if(_stream_matmul_55_stream_oready) begin
        _tmp_1932 <= _stream_matmul_55_sink_busy;
      end 
      if(!_stream_matmul_55_sink_busy && _tmp_1932) begin
        _stream_matmul_55_busy_reg <= 0;
      end 
      if(_stream_matmul_55_source_busy) begin
        _stream_matmul_55_busy_reg <= 1;
      end 
    end
  end

  localparam _stream_matmul_55_fsm_1 = 1;
  localparam _stream_matmul_55_fsm_2 = 2;
  localparam _stream_matmul_55_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_matmul_55_fsm <= _stream_matmul_55_fsm_init;
      _stream_matmul_55_source_start <= 0;
      _stream_matmul_55_source_busy <= 0;
      _stream_matmul_55_stream_ivalid <= 0;
    end else begin
      if(_stream_matmul_55_stream_oready && _tmp_1825) begin
        _stream_matmul_55_stream_ivalid <= 1;
      end 
      if(_stream_matmul_55_stream_oready && _tmp_1835) begin
        _stream_matmul_55_stream_ivalid <= 0;
      end 
      case(_stream_matmul_55_fsm)
        _stream_matmul_55_fsm_init: begin
          if(_stream_matmul_55_run_flag) begin
            _stream_matmul_55_source_start <= 1;
          end 
          if(_stream_matmul_55_run_flag) begin
            _stream_matmul_55_fsm <= _stream_matmul_55_fsm_1;
          end 
        end
        _stream_matmul_55_fsm_1: begin
          if(_stream_matmul_55_source_start && _stream_matmul_55_stream_oready) begin
            _stream_matmul_55_source_start <= 0;
            _stream_matmul_55_source_busy <= 1;
          end 
          if(_stream_matmul_55_source_start && _stream_matmul_55_stream_oready) begin
            _stream_matmul_55_fsm <= _stream_matmul_55_fsm_2;
          end 
        end
        _stream_matmul_55_fsm_2: begin
          if(_stream_matmul_55_stream_oready) begin
            _stream_matmul_55_fsm <= _stream_matmul_55_fsm_3;
          end 
        end
        _stream_matmul_55_fsm_3: begin
          if(_stream_matmul_55_stream_oready && (_stream_matmul_55_source_11_idle && _stream_matmul_55_source_13_idle && _stream_matmul_55_source_15_idle && _stream_matmul_55_source_20_idle && _stream_matmul_55_source_21_idle && _stream_matmul_55_source_7_idle && _stream_matmul_55_source_9_idle && (_stream_matmul_55_fsm == 3))) begin
            _stream_matmul_55_source_busy <= 0;
          end 
          if(_stream_matmul_55_stream_oready && (_stream_matmul_55_source_11_idle && _stream_matmul_55_source_13_idle && _stream_matmul_55_source_15_idle && _stream_matmul_55_source_20_idle && _stream_matmul_55_source_21_idle && _stream_matmul_55_source_7_idle && _stream_matmul_55_source_9_idle && (_stream_matmul_55_fsm == 3)) && _stream_matmul_55_run_flag) begin
            _stream_matmul_55_source_start <= 1;
          end 
          if(_stream_matmul_55_stream_oready && (_stream_matmul_55_source_11_idle && _stream_matmul_55_source_13_idle && _stream_matmul_55_source_15_idle && _stream_matmul_55_source_20_idle && _stream_matmul_55_source_21_idle && _stream_matmul_55_source_7_idle && _stream_matmul_55_source_9_idle && (_stream_matmul_55_fsm == 3))) begin
            _stream_matmul_55_fsm <= _stream_matmul_55_fsm_init;
          end 
          if(_stream_matmul_55_stream_oready && (_stream_matmul_55_source_11_idle && _stream_matmul_55_source_13_idle && _stream_matmul_55_source_15_idle && _stream_matmul_55_source_20_idle && _stream_matmul_55_source_21_idle && _stream_matmul_55_source_7_idle && _stream_matmul_55_source_9_idle && (_stream_matmul_55_fsm == 3)) && _stream_matmul_55_run_flag) begin
            _stream_matmul_55_fsm <= _stream_matmul_55_fsm_1;
          end 
        end
      endcase
    end
  end

  localparam main_fsm_1 = 1;
  localparam main_fsm_2 = 2;
  localparam main_fsm_3 = 3;
  localparam main_fsm_4 = 4;
  localparam main_fsm_5 = 5;
  localparam main_fsm_6 = 6;
  localparam main_fsm_7 = 7;
  localparam main_fsm_8 = 8;
  localparam main_fsm_9 = 9;
  localparam main_fsm_10 = 10;
  localparam main_fsm_11 = 11;
  localparam main_fsm_12 = 12;
  localparam main_fsm_13 = 13;
  localparam main_fsm_14 = 14;
  localparam main_fsm_15 = 15;
  localparam main_fsm_16 = 16;
  localparam main_fsm_17 = 17;
  localparam main_fsm_18 = 18;
  localparam main_fsm_19 = 19;
  localparam main_fsm_20 = 20;
  localparam main_fsm_21 = 21;
  localparam main_fsm_22 = 22;
  localparam main_fsm_23 = 23;
  localparam main_fsm_24 = 24;
  localparam main_fsm_25 = 25;
  localparam main_fsm_26 = 26;
  localparam main_fsm_27 = 27;
  localparam main_fsm_28 = 28;
  localparam main_fsm_29 = 29;
  localparam main_fsm_30 = 30;
  localparam main_fsm_31 = 31;
  localparam main_fsm_32 = 32;
  localparam main_fsm_33 = 33;
  localparam main_fsm_34 = 34;
  localparam main_fsm_35 = 35;
  localparam main_fsm_36 = 36;
  localparam main_fsm_37 = 37;
  localparam main_fsm_38 = 38;
  localparam main_fsm_39 = 39;
  localparam main_fsm_40 = 40;
  localparam main_fsm_41 = 41;
  localparam main_fsm_42 = 42;
  localparam main_fsm_43 = 43;
  localparam main_fsm_44 = 44;
  localparam main_fsm_45 = 45;
  localparam main_fsm_46 = 46;
  localparam main_fsm_47 = 47;
  localparam main_fsm_48 = 48;
  localparam main_fsm_49 = 49;
  localparam main_fsm_50 = 50;
  localparam main_fsm_51 = 51;
  localparam main_fsm_52 = 52;
  localparam main_fsm_53 = 53;
  localparam main_fsm_54 = 54;
  localparam main_fsm_55 = 55;
  localparam main_fsm_56 = 56;
  localparam main_fsm_57 = 57;
  localparam main_fsm_58 = 58;
  localparam main_fsm_59 = 59;
  localparam main_fsm_60 = 60;
  localparam main_fsm_61 = 61;
  localparam main_fsm_62 = 62;
  localparam main_fsm_63 = 63;
  localparam main_fsm_64 = 64;
  localparam main_fsm_65 = 65;
  localparam main_fsm_66 = 66;
  localparam main_fsm_67 = 67;
  localparam main_fsm_68 = 68;
  localparam main_fsm_69 = 69;
  localparam main_fsm_70 = 70;
  localparam main_fsm_71 = 71;
  localparam main_fsm_72 = 72;
  localparam main_fsm_73 = 73;
  localparam main_fsm_74 = 74;
  localparam main_fsm_75 = 75;
  localparam main_fsm_76 = 76;
  localparam main_fsm_77 = 77;
  localparam main_fsm_78 = 78;
  localparam main_fsm_79 = 79;
  localparam main_fsm_80 = 80;
  localparam main_fsm_81 = 81;
  localparam main_fsm_82 = 82;
  localparam main_fsm_83 = 83;
  localparam main_fsm_84 = 84;
  localparam main_fsm_85 = 85;
  localparam main_fsm_86 = 86;
  localparam main_fsm_87 = 87;
  localparam main_fsm_88 = 88;
  localparam main_fsm_89 = 89;
  localparam main_fsm_90 = 90;
  localparam main_fsm_91 = 91;
  localparam main_fsm_92 = 92;
  localparam main_fsm_93 = 93;
  localparam main_fsm_94 = 94;
  localparam main_fsm_95 = 95;
  localparam main_fsm_96 = 96;
  localparam main_fsm_97 = 97;
  localparam main_fsm_98 = 98;
  localparam main_fsm_99 = 99;
  localparam main_fsm_100 = 100;
  localparam main_fsm_101 = 101;
  localparam main_fsm_102 = 102;
  localparam main_fsm_103 = 103;
  localparam main_fsm_104 = 104;
  localparam main_fsm_105 = 105;
  localparam main_fsm_106 = 106;
  localparam main_fsm_107 = 107;
  localparam main_fsm_108 = 108;
  localparam main_fsm_109 = 109;
  localparam main_fsm_110 = 110;
  localparam main_fsm_111 = 111;
  localparam main_fsm_112 = 112;
  localparam main_fsm_113 = 113;
  localparam main_fsm_114 = 114;
  localparam main_fsm_115 = 115;
  localparam main_fsm_116 = 116;
  localparam main_fsm_117 = 117;
  localparam main_fsm_118 = 118;
  localparam main_fsm_119 = 119;
  localparam main_fsm_120 = 120;
  localparam main_fsm_121 = 121;
  localparam main_fsm_122 = 122;
  localparam main_fsm_123 = 123;
  localparam main_fsm_124 = 124;
  localparam main_fsm_125 = 125;
  localparam main_fsm_126 = 126;
  localparam main_fsm_127 = 127;
  localparam main_fsm_128 = 128;
  localparam main_fsm_129 = 129;
  localparam main_fsm_130 = 130;
  localparam main_fsm_131 = 131;
  localparam main_fsm_132 = 132;
  localparam main_fsm_133 = 133;
  localparam main_fsm_134 = 134;
  localparam main_fsm_135 = 135;
  localparam main_fsm_136 = 136;
  localparam main_fsm_137 = 137;
  localparam main_fsm_138 = 138;
  localparam main_fsm_139 = 139;
  localparam main_fsm_140 = 140;
  localparam main_fsm_141 = 141;
  localparam main_fsm_142 = 142;
  localparam main_fsm_143 = 143;
  localparam main_fsm_144 = 144;
  localparam main_fsm_145 = 145;
  localparam main_fsm_146 = 146;
  localparam main_fsm_147 = 147;
  localparam main_fsm_148 = 148;
  localparam main_fsm_149 = 149;
  localparam main_fsm_150 = 150;
  localparam main_fsm_151 = 151;
  localparam main_fsm_152 = 152;
  localparam main_fsm_153 = 153;
  localparam main_fsm_154 = 154;
  localparam main_fsm_155 = 155;
  localparam main_fsm_156 = 156;
  localparam main_fsm_157 = 157;
  localparam main_fsm_158 = 158;
  localparam main_fsm_159 = 159;
  localparam main_fsm_160 = 160;
  localparam main_fsm_161 = 161;
  localparam main_fsm_162 = 162;

  always @(posedge CLK) begin
    if(RST) begin
      main_fsm <= main_fsm_init;
      conv2d_24_objaddr <= 0;
      conv2d_24_arg_objaddr_0 <= 0;
      conv2d_24_arg_objaddr_1 <= 0;
      conv2d_24_arg_objaddr_2 <= 0;
      conv2d_24_arg_objaddr_3 <= 0;
      conv2d_24_control_param_index <= 0;
      max_pool_serial_26_objaddr <= 0;
      max_pool_serial_26_arg_objaddr_0 <= 0;
      max_pool_serial_26_control_param_index <= 0;
      avg_pool_serial_52_objaddr <= 0;
      avg_pool_serial_52_arg_objaddr_0 <= 0;
      matmul_55_objaddr <= 0;
      matmul_55_arg_objaddr_0 <= 0;
      matmul_55_arg_objaddr_1 <= 0;
      matmul_55_arg_objaddr_2 <= 0;
      matmul_55_arg_objaddr_3 <= 0;
      matmul_55_control_param_index <= 0;
    end else begin
      case(main_fsm)
        main_fsm_init: begin
          if(_saxi_register_4 != 0) begin
            main_fsm <= main_fsm_1;
          end 
        end
        main_fsm_1: begin
          main_fsm <= main_fsm_2;
        end
        main_fsm_2: begin
          main_fsm <= main_fsm_3;
        end
        main_fsm_3: begin
          main_fsm <= main_fsm_4;
        end
        main_fsm_4: begin
          main_fsm <= main_fsm_5;
        end
        main_fsm_5: begin
          conv2d_24_objaddr <= _saxi_register_33;
          main_fsm <= main_fsm_6;
        end
        main_fsm_6: begin
          conv2d_24_arg_objaddr_0 <= _saxi_register_35;
          main_fsm <= main_fsm_7;
        end
        main_fsm_7: begin
          conv2d_24_arg_objaddr_1 <= _saxi_register_36;
          main_fsm <= main_fsm_8;
        end
        main_fsm_8: begin
          conv2d_24_arg_objaddr_2 <= _saxi_register_36 + 2304;
          main_fsm <= main_fsm_9;
        end
        main_fsm_9: begin
          conv2d_24_arg_objaddr_3 <= _saxi_register_36 + 2560;
          main_fsm <= main_fsm_10;
        end
        main_fsm_10: begin
          conv2d_24_control_param_index <= 0;
          main_fsm <= main_fsm_11;
        end
        main_fsm_11: begin
          main_fsm <= main_fsm_12;
        end
        main_fsm_12: begin
          main_fsm <= main_fsm_13;
        end
        main_fsm_13: begin
          if(control_conv2d_24 == 34) begin
            main_fsm <= main_fsm_14;
          end 
        end
        main_fsm_14: begin
          main_fsm <= main_fsm_15;
        end
        main_fsm_15: begin
          max_pool_serial_26_objaddr <= _saxi_register_33 + 3211264;
          main_fsm <= main_fsm_16;
        end
        main_fsm_16: begin
          max_pool_serial_26_arg_objaddr_0 <= _saxi_register_33;
          main_fsm <= main_fsm_17;
        end
        main_fsm_17: begin
          max_pool_serial_26_control_param_index <= 0;
          main_fsm <= main_fsm_18;
        end
        main_fsm_18: begin
          main_fsm <= main_fsm_19;
        end
        main_fsm_19: begin
          main_fsm <= main_fsm_20;
        end
        main_fsm_20: begin
          if(control_max_pool_serial_26 == 19) begin
            main_fsm <= main_fsm_21;
          end 
        end
        main_fsm_21: begin
          main_fsm <= main_fsm_22;
        end
        main_fsm_22: begin
          conv2d_24_objaddr <= _saxi_register_33 + 4014080;
          main_fsm <= main_fsm_23;
        end
        main_fsm_23: begin
          conv2d_24_arg_objaddr_0 <= _saxi_register_33 + 3211264;
          main_fsm <= main_fsm_24;
        end
        main_fsm_24: begin
          conv2d_24_arg_objaddr_1 <= _saxi_register_36 + 2624;
          main_fsm <= main_fsm_25;
        end
        main_fsm_25: begin
          conv2d_24_arg_objaddr_2 <= _saxi_register_36 + 76352;
          main_fsm <= main_fsm_26;
        end
        main_fsm_26: begin
          conv2d_24_arg_objaddr_3 <= _saxi_register_36 + 76864;
          main_fsm <= main_fsm_27;
        end
        main_fsm_27: begin
          conv2d_24_control_param_index <= 1;
          main_fsm <= main_fsm_28;
        end
        main_fsm_28: begin
          main_fsm <= main_fsm_29;
        end
        main_fsm_29: begin
          main_fsm <= main_fsm_30;
        end
        main_fsm_30: begin
          if(control_conv2d_24 == 34) begin
            main_fsm <= main_fsm_31;
          end 
        end
        main_fsm_31: begin
          main_fsm <= main_fsm_32;
        end
        main_fsm_32: begin
          max_pool_serial_26_objaddr <= _saxi_register_33 + 5619712;
          main_fsm <= main_fsm_33;
        end
        main_fsm_33: begin
          max_pool_serial_26_arg_objaddr_0 <= _saxi_register_33 + 4014080;
          main_fsm <= main_fsm_34;
        end
        main_fsm_34: begin
          max_pool_serial_26_control_param_index <= 1;
          main_fsm <= main_fsm_35;
        end
        main_fsm_35: begin
          main_fsm <= main_fsm_36;
        end
        main_fsm_36: begin
          main_fsm <= main_fsm_37;
        end
        main_fsm_37: begin
          if(control_max_pool_serial_26 == 19) begin
            main_fsm <= main_fsm_38;
          end 
        end
        main_fsm_38: begin
          main_fsm <= main_fsm_39;
        end
        main_fsm_39: begin
          conv2d_24_objaddr <= _saxi_register_33 + 6021120;
          main_fsm <= main_fsm_40;
        end
        main_fsm_40: begin
          conv2d_24_arg_objaddr_0 <= _saxi_register_33 + 5619712;
          main_fsm <= main_fsm_41;
        end
        main_fsm_41: begin
          conv2d_24_arg_objaddr_1 <= _saxi_register_36 + 76928;
          main_fsm <= main_fsm_42;
        end
        main_fsm_42: begin
          conv2d_24_arg_objaddr_2 <= _saxi_register_36 + 371840;
          main_fsm <= main_fsm_43;
        end
        main_fsm_43: begin
          conv2d_24_arg_objaddr_3 <= _saxi_register_36 + 372864;
          main_fsm <= main_fsm_44;
        end
        main_fsm_44: begin
          conv2d_24_control_param_index <= 2;
          main_fsm <= main_fsm_45;
        end
        main_fsm_45: begin
          main_fsm <= main_fsm_46;
        end
        main_fsm_46: begin
          main_fsm <= main_fsm_47;
        end
        main_fsm_47: begin
          if(control_conv2d_24 == 34) begin
            main_fsm <= main_fsm_48;
          end 
        end
        main_fsm_48: begin
          main_fsm <= main_fsm_49;
        end
        main_fsm_49: begin
          conv2d_24_objaddr <= _saxi_register_33 + 6823936;
          main_fsm <= main_fsm_50;
        end
        main_fsm_50: begin
          conv2d_24_arg_objaddr_0 <= _saxi_register_33 + 6021120;
          main_fsm <= main_fsm_51;
        end
        main_fsm_51: begin
          conv2d_24_arg_objaddr_1 <= _saxi_register_36 + 372928;
          main_fsm <= main_fsm_52;
        end
        main_fsm_52: begin
          conv2d_24_arg_objaddr_2 <= _saxi_register_36 + 962752;
          main_fsm <= main_fsm_53;
        end
        main_fsm_53: begin
          conv2d_24_arg_objaddr_3 <= _saxi_register_36 + 963776;
          main_fsm <= main_fsm_54;
        end
        main_fsm_54: begin
          conv2d_24_control_param_index <= 3;
          main_fsm <= main_fsm_55;
        end
        main_fsm_55: begin
          main_fsm <= main_fsm_56;
        end
        main_fsm_56: begin
          main_fsm <= main_fsm_57;
        end
        main_fsm_57: begin
          if(control_conv2d_24 == 34) begin
            main_fsm <= main_fsm_58;
          end 
        end
        main_fsm_58: begin
          main_fsm <= main_fsm_59;
        end
        main_fsm_59: begin
          max_pool_serial_26_objaddr <= _saxi_register_33 + 7626752;
          main_fsm <= main_fsm_60;
        end
        main_fsm_60: begin
          max_pool_serial_26_arg_objaddr_0 <= _saxi_register_33 + 6823936;
          main_fsm <= main_fsm_61;
        end
        main_fsm_61: begin
          max_pool_serial_26_control_param_index <= 2;
          main_fsm <= main_fsm_62;
        end
        main_fsm_62: begin
          main_fsm <= main_fsm_63;
        end
        main_fsm_63: begin
          main_fsm <= main_fsm_64;
        end
        main_fsm_64: begin
          if(control_max_pool_serial_26 == 19) begin
            main_fsm <= main_fsm_65;
          end 
        end
        main_fsm_65: begin
          main_fsm <= main_fsm_66;
        end
        main_fsm_66: begin
          conv2d_24_objaddr <= _saxi_register_33 + 7827456;
          main_fsm <= main_fsm_67;
        end
        main_fsm_67: begin
          conv2d_24_arg_objaddr_0 <= _saxi_register_33 + 7626752;
          main_fsm <= main_fsm_68;
        end
        main_fsm_68: begin
          conv2d_24_arg_objaddr_1 <= _saxi_register_36 + 963840;
          main_fsm <= main_fsm_69;
        end
        main_fsm_69: begin
          conv2d_24_arg_objaddr_2 <= _saxi_register_36 + 2143488;
          main_fsm <= main_fsm_70;
        end
        main_fsm_70: begin
          conv2d_24_arg_objaddr_3 <= _saxi_register_36 + 2145536;
          main_fsm <= main_fsm_71;
        end
        main_fsm_71: begin
          conv2d_24_control_param_index <= 4;
          main_fsm <= main_fsm_72;
        end
        main_fsm_72: begin
          main_fsm <= main_fsm_73;
        end
        main_fsm_73: begin
          main_fsm <= main_fsm_74;
        end
        main_fsm_74: begin
          if(control_conv2d_24 == 34) begin
            main_fsm <= main_fsm_75;
          end 
        end
        main_fsm_75: begin
          main_fsm <= main_fsm_76;
        end
        main_fsm_76: begin
          conv2d_24_objaddr <= _saxi_register_33 + 8228864;
          main_fsm <= main_fsm_77;
        end
        main_fsm_77: begin
          conv2d_24_arg_objaddr_0 <= _saxi_register_33 + 7827456;
          main_fsm <= main_fsm_78;
        end
        main_fsm_78: begin
          conv2d_24_arg_objaddr_1 <= _saxi_register_36 + 2145600;
          main_fsm <= main_fsm_79;
        end
        main_fsm_79: begin
          conv2d_24_arg_objaddr_2 <= _saxi_register_36 + 4504896;
          main_fsm <= main_fsm_80;
        end
        main_fsm_80: begin
          conv2d_24_arg_objaddr_3 <= _saxi_register_36 + 4506944;
          main_fsm <= main_fsm_81;
        end
        main_fsm_81: begin
          conv2d_24_control_param_index <= 5;
          main_fsm <= main_fsm_82;
        end
        main_fsm_82: begin
          main_fsm <= main_fsm_83;
        end
        main_fsm_83: begin
          main_fsm <= main_fsm_84;
        end
        main_fsm_84: begin
          if(control_conv2d_24 == 34) begin
            main_fsm <= main_fsm_85;
          end 
        end
        main_fsm_85: begin
          main_fsm <= main_fsm_86;
        end
        main_fsm_86: begin
          max_pool_serial_26_objaddr <= _saxi_register_33 + 8630272;
          main_fsm <= main_fsm_87;
        end
        main_fsm_87: begin
          max_pool_serial_26_arg_objaddr_0 <= _saxi_register_33 + 8228864;
          main_fsm <= main_fsm_88;
        end
        main_fsm_88: begin
          max_pool_serial_26_control_param_index <= 3;
          main_fsm <= main_fsm_89;
        end
        main_fsm_89: begin
          main_fsm <= main_fsm_90;
        end
        main_fsm_90: begin
          main_fsm <= main_fsm_91;
        end
        main_fsm_91: begin
          if(control_max_pool_serial_26 == 19) begin
            main_fsm <= main_fsm_92;
          end 
        end
        main_fsm_92: begin
          main_fsm <= main_fsm_93;
        end
        main_fsm_93: begin
          conv2d_24_objaddr <= _saxi_register_33 + 8730624;
          main_fsm <= main_fsm_94;
        end
        main_fsm_94: begin
          conv2d_24_arg_objaddr_0 <= _saxi_register_33 + 8630272;
          main_fsm <= main_fsm_95;
        end
        main_fsm_95: begin
          conv2d_24_arg_objaddr_1 <= _saxi_register_36 + 4507008;
          main_fsm <= main_fsm_96;
        end
        main_fsm_96: begin
          conv2d_24_arg_objaddr_2 <= _saxi_register_36 + 6866304;
          main_fsm <= main_fsm_97;
        end
        main_fsm_97: begin
          conv2d_24_arg_objaddr_3 <= _saxi_register_36 + 6868352;
          main_fsm <= main_fsm_98;
        end
        main_fsm_98: begin
          conv2d_24_control_param_index <= 6;
          main_fsm <= main_fsm_99;
        end
        main_fsm_99: begin
          main_fsm <= main_fsm_100;
        end
        main_fsm_100: begin
          main_fsm <= main_fsm_101;
        end
        main_fsm_101: begin
          if(control_conv2d_24 == 34) begin
            main_fsm <= main_fsm_102;
          end 
        end
        main_fsm_102: begin
          main_fsm <= main_fsm_103;
        end
        main_fsm_103: begin
          conv2d_24_objaddr <= _saxi_register_33 + 8830976;
          main_fsm <= main_fsm_104;
        end
        main_fsm_104: begin
          conv2d_24_arg_objaddr_0 <= _saxi_register_33 + 8730624;
          main_fsm <= main_fsm_105;
        end
        main_fsm_105: begin
          conv2d_24_arg_objaddr_1 <= _saxi_register_36 + 6868416;
          main_fsm <= main_fsm_106;
        end
        main_fsm_106: begin
          conv2d_24_arg_objaddr_2 <= _saxi_register_36 + 9227712;
          main_fsm <= main_fsm_107;
        end
        main_fsm_107: begin
          conv2d_24_arg_objaddr_3 <= _saxi_register_36 + 9229760;
          main_fsm <= main_fsm_108;
        end
        main_fsm_108: begin
          conv2d_24_control_param_index <= 7;
          main_fsm <= main_fsm_109;
        end
        main_fsm_109: begin
          main_fsm <= main_fsm_110;
        end
        main_fsm_110: begin
          main_fsm <= main_fsm_111;
        end
        main_fsm_111: begin
          if(control_conv2d_24 == 34) begin
            main_fsm <= main_fsm_112;
          end 
        end
        main_fsm_112: begin
          main_fsm <= main_fsm_113;
        end
        main_fsm_113: begin
          max_pool_serial_26_objaddr <= _saxi_register_33 + 8931328;
          main_fsm <= main_fsm_114;
        end
        main_fsm_114: begin
          max_pool_serial_26_arg_objaddr_0 <= _saxi_register_33 + 8830976;
          main_fsm <= main_fsm_115;
        end
        main_fsm_115: begin
          max_pool_serial_26_control_param_index <= 4;
          main_fsm <= main_fsm_116;
        end
        main_fsm_116: begin
          main_fsm <= main_fsm_117;
        end
        main_fsm_117: begin
          main_fsm <= main_fsm_118;
        end
        main_fsm_118: begin
          if(control_max_pool_serial_26 == 19) begin
            main_fsm <= main_fsm_119;
          end 
        end
        main_fsm_119: begin
          main_fsm <= main_fsm_120;
        end
        main_fsm_120: begin
          avg_pool_serial_52_objaddr <= _saxi_register_33 + 8956416;
          main_fsm <= main_fsm_121;
        end
        main_fsm_121: begin
          avg_pool_serial_52_arg_objaddr_0 <= _saxi_register_33 + 8931328;
          main_fsm <= main_fsm_122;
        end
        main_fsm_122: begin
          main_fsm <= main_fsm_123;
        end
        main_fsm_123: begin
          main_fsm <= main_fsm_124;
        end
        main_fsm_124: begin
          if(control_avg_pool_serial_52 == 16) begin
            main_fsm <= main_fsm_125;
          end 
        end
        main_fsm_125: begin
          main_fsm <= main_fsm_126;
        end
        main_fsm_126: begin
          main_fsm <= main_fsm_127;
        end
        main_fsm_127: begin
          main_fsm <= main_fsm_128;
        end
        main_fsm_128: begin
          matmul_55_objaddr <= _saxi_register_33 + 8981504;
          main_fsm <= main_fsm_129;
        end
        main_fsm_129: begin
          matmul_55_arg_objaddr_0 <= _saxi_register_33 + 8956416;
          main_fsm <= main_fsm_130;
        end
        main_fsm_130: begin
          matmul_55_arg_objaddr_1 <= _saxi_register_36 + 9229824;
          main_fsm <= main_fsm_131;
        end
        main_fsm_131: begin
          matmul_55_arg_objaddr_2 <= _saxi_register_36 + 111990272;
          main_fsm <= main_fsm_132;
        end
        main_fsm_132: begin
          matmul_55_arg_objaddr_3 <= _saxi_register_36 + 112006656;
          main_fsm <= main_fsm_133;
        end
        main_fsm_133: begin
          matmul_55_control_param_index <= 0;
          main_fsm <= main_fsm_134;
        end
        main_fsm_134: begin
          main_fsm <= main_fsm_135;
        end
        main_fsm_135: begin
          main_fsm <= main_fsm_136;
        end
        main_fsm_136: begin
          if(control_matmul_55 == 28) begin
            main_fsm <= main_fsm_137;
          end 
        end
        main_fsm_137: begin
          main_fsm <= main_fsm_138;
        end
        main_fsm_138: begin
          matmul_55_objaddr <= _saxi_register_33 + 8985600;
          main_fsm <= main_fsm_139;
        end
        main_fsm_139: begin
          matmul_55_arg_objaddr_0 <= _saxi_register_33 + 8981504;
          main_fsm <= main_fsm_140;
        end
        main_fsm_140: begin
          matmul_55_arg_objaddr_1 <= _saxi_register_36 + 112006720;
          main_fsm <= main_fsm_141;
        end
        main_fsm_141: begin
          matmul_55_arg_objaddr_2 <= _saxi_register_36 + 128783936;
          main_fsm <= main_fsm_142;
        end
        main_fsm_142: begin
          matmul_55_arg_objaddr_3 <= _saxi_register_36 + 128800320;
          main_fsm <= main_fsm_143;
        end
        main_fsm_143: begin
          matmul_55_control_param_index <= 1;
          main_fsm <= main_fsm_144;
        end
        main_fsm_144: begin
          main_fsm <= main_fsm_145;
        end
        main_fsm_145: begin
          main_fsm <= main_fsm_146;
        end
        main_fsm_146: begin
          if(control_matmul_55 == 28) begin
            main_fsm <= main_fsm_147;
          end 
        end
        main_fsm_147: begin
          main_fsm <= main_fsm_148;
        end
        main_fsm_148: begin
          matmul_55_objaddr <= _saxi_register_34;
          main_fsm <= main_fsm_149;
        end
        main_fsm_149: begin
          matmul_55_arg_objaddr_0 <= _saxi_register_33 + 8985600;
          main_fsm <= main_fsm_150;
        end
        main_fsm_150: begin
          matmul_55_arg_objaddr_1 <= _saxi_register_36 + 128800384;
          main_fsm <= main_fsm_151;
        end
        main_fsm_151: begin
          matmul_55_arg_objaddr_2 <= _saxi_register_36 + 132896384;
          main_fsm <= main_fsm_152;
        end
        main_fsm_152: begin
          matmul_55_arg_objaddr_3 <= _saxi_register_36 + 132900416;
          main_fsm <= main_fsm_153;
        end
        main_fsm_153: begin
          matmul_55_control_param_index <= 2;
          main_fsm <= main_fsm_154;
        end
        main_fsm_154: begin
          main_fsm <= main_fsm_155;
        end
        main_fsm_155: begin
          main_fsm <= main_fsm_156;
        end
        main_fsm_156: begin
          if(control_matmul_55 == 28) begin
            main_fsm <= main_fsm_157;
          end 
        end
        main_fsm_157: begin
          main_fsm <= main_fsm_158;
        end
        main_fsm_158: begin
          main_fsm <= main_fsm_159;
        end
        main_fsm_159: begin
          main_fsm <= main_fsm_160;
        end
        main_fsm_160: begin
          main_fsm <= main_fsm_161;
        end
        main_fsm_161: begin
          main_fsm <= main_fsm_162;
        end
        main_fsm_162: begin
          main_fsm <= main_fsm_init;
        end
      endcase
    end
  end

  localparam control_conv2d_24_1 = 1;
  localparam control_conv2d_24_2 = 2;
  localparam control_conv2d_24_3 = 3;
  localparam control_conv2d_24_4 = 4;
  localparam control_conv2d_24_5 = 5;
  localparam control_conv2d_24_6 = 6;
  localparam control_conv2d_24_7 = 7;
  localparam control_conv2d_24_8 = 8;
  localparam control_conv2d_24_9 = 9;
  localparam control_conv2d_24_10 = 10;
  localparam control_conv2d_24_11 = 11;
  localparam control_conv2d_24_12 = 12;
  localparam control_conv2d_24_13 = 13;
  localparam control_conv2d_24_14 = 14;
  localparam control_conv2d_24_15 = 15;
  localparam control_conv2d_24_16 = 16;
  localparam control_conv2d_24_17 = 17;
  localparam control_conv2d_24_18 = 18;
  localparam control_conv2d_24_19 = 19;
  localparam control_conv2d_24_20 = 20;
  localparam control_conv2d_24_21 = 21;
  localparam control_conv2d_24_22 = 22;
  localparam control_conv2d_24_23 = 23;
  localparam control_conv2d_24_24 = 24;
  localparam control_conv2d_24_25 = 25;
  localparam control_conv2d_24_26 = 26;
  localparam control_conv2d_24_27 = 27;
  localparam control_conv2d_24_28 = 28;
  localparam control_conv2d_24_29 = 29;
  localparam control_conv2d_24_30 = 30;
  localparam control_conv2d_24_31 = 31;
  localparam control_conv2d_24_32 = 32;
  localparam control_conv2d_24_33 = 33;
  localparam control_conv2d_24_34 = 34;

  always @(posedge CLK) begin
    if(RST) begin
      control_conv2d_24 <= control_conv2d_24_init;
      _control_conv2d_24_called <= 0;
      conv2d_24_filter_base_offset <= 0;
      conv2d_24_filter_page_comp_offset <= 0;
      conv2d_24_filter_page_dma_offset <= 0;
      conv2d_24_act_base_offset_row <= 0;
      conv2d_24_act_base_offset_bat <= 0;
      conv2d_24_dma_flag_0 <= 0;
      conv2d_24_dma_flag_1 <= 0;
      conv2d_24_dma_flag_2 <= 0;
      conv2d_24_act_page_comp_offset_0 <= 0;
      conv2d_24_act_page_comp_offset_1 <= 0;
      conv2d_24_act_page_comp_offset_2 <= 0;
      conv2d_24_act_page_dma_offset_0 <= 0;
      conv2d_24_act_page_dma_offset_1 <= 0;
      conv2d_24_act_page_dma_offset_2 <= 0;
      conv2d_24_out_base_offset_val <= 0;
      conv2d_24_out_base_offset_col <= 0;
      conv2d_24_out_base_offset_row <= 0;
      conv2d_24_out_base_offset_bat <= 0;
      conv2d_24_out_base_offset_och <= 0;
      conv2d_24_out_page <= 0;
      conv2d_24_out_page_comp_offset <= 0;
      conv2d_24_out_page_dma_offset <= 0;
      conv2d_24_out_laddr_offset <= 0;
      conv2d_24_sync_out_count <= 0;
      conv2d_24_write_count <= 0;
      conv2d_24_next_out_write_size <= 0;
      conv2d_24_row_count <= 0;
      conv2d_24_bat_count <= 0;
      conv2d_24_och_count <= 0;
      conv2d_24_row_select <= 0;
      conv2d_24_prev_row_count <= 0;
      conv2d_24_prev_bat_count <= 0;
      conv2d_24_prev_och_count <= 0;
      conv2d_24_prev_row_select <= 0;
      conv2d_24_out_col_count <= 0;
      conv2d_24_out_row_count <= 0;
      conv2d_24_out_ram_select <= 0;
      conv2d_24_skip_read_filter <= 0;
      conv2d_24_skip_read_act <= 0;
      conv2d_24_skip_comp <= 0;
      conv2d_24_skip_write_out <= 1;
    end else begin
      case(control_conv2d_24)
        control_conv2d_24_init: begin
          if(main_fsm == 11) begin
            _control_conv2d_24_called <= 1;
          end 
          if(main_fsm == 28) begin
            _control_conv2d_24_called <= 1;
          end 
          if(main_fsm == 45) begin
            _control_conv2d_24_called <= 1;
          end 
          if(main_fsm == 55) begin
            _control_conv2d_24_called <= 1;
          end 
          if(main_fsm == 72) begin
            _control_conv2d_24_called <= 1;
          end 
          if(main_fsm == 82) begin
            _control_conv2d_24_called <= 1;
          end 
          if(main_fsm == 99) begin
            _control_conv2d_24_called <= 1;
          end 
          if(main_fsm == 109) begin
            _control_conv2d_24_called <= 1;
          end 
          if(main_fsm == 11) begin
            control_conv2d_24 <= control_conv2d_24_1;
          end 
          if(main_fsm == 28) begin
            control_conv2d_24 <= control_conv2d_24_1;
          end 
          if(main_fsm == 45) begin
            control_conv2d_24 <= control_conv2d_24_1;
          end 
          if(main_fsm == 55) begin
            control_conv2d_24 <= control_conv2d_24_1;
          end 
          if(main_fsm == 72) begin
            control_conv2d_24 <= control_conv2d_24_1;
          end 
          if(main_fsm == 82) begin
            control_conv2d_24 <= control_conv2d_24_1;
          end 
          if(main_fsm == 99) begin
            control_conv2d_24 <= control_conv2d_24_1;
          end 
          if(main_fsm == 109) begin
            control_conv2d_24 <= control_conv2d_24_1;
          end 
        end
        control_conv2d_24_1: begin
          control_conv2d_24 <= control_conv2d_24_2;
        end
        control_conv2d_24_2: begin
          conv2d_24_filter_base_offset <= 0;
          conv2d_24_filter_page_comp_offset <= 0;
          conv2d_24_filter_page_dma_offset <= 0;
          conv2d_24_act_base_offset_row <= 0;
          conv2d_24_act_base_offset_bat <= 0;
          conv2d_24_dma_flag_0 <= 1;
          conv2d_24_dma_flag_1 <= 1;
          conv2d_24_dma_flag_2 <= 1;
          conv2d_24_act_page_comp_offset_0 <= 0;
          conv2d_24_act_page_comp_offset_1 <= 0;
          conv2d_24_act_page_comp_offset_2 <= 0;
          conv2d_24_act_page_dma_offset_0 <= 0;
          conv2d_24_act_page_dma_offset_1 <= 0;
          conv2d_24_act_page_dma_offset_2 <= 0;
          conv2d_24_out_base_offset_val <= 0;
          conv2d_24_out_base_offset_col <= 0;
          conv2d_24_out_base_offset_row <= 0;
          conv2d_24_out_base_offset_bat <= 0;
          conv2d_24_out_base_offset_och <= 0;
          conv2d_24_out_page <= 0;
          conv2d_24_out_page_comp_offset <= 0;
          conv2d_24_out_page_dma_offset <= 0;
          conv2d_24_out_laddr_offset <= 0;
          conv2d_24_sync_out_count <= 0;
          conv2d_24_write_count <= 0;
          conv2d_24_next_out_write_size <= (cparam_conv2d_24_max_och_count == 0)? cparam_conv2d_24_out_write_size_res : cparam_conv2d_24_out_write_size;
          conv2d_24_row_count <= 0;
          conv2d_24_bat_count <= 0;
          conv2d_24_och_count <= 0;
          conv2d_24_row_select <= 0;
          conv2d_24_prev_row_count <= 0;
          conv2d_24_prev_bat_count <= 0;
          conv2d_24_prev_och_count <= 0;
          conv2d_24_prev_row_select <= 0;
          conv2d_24_out_col_count <= 0;
          conv2d_24_out_row_count <= 0;
          conv2d_24_out_ram_select <= 0;
          conv2d_24_skip_read_filter <= 0;
          conv2d_24_skip_read_act <= 0;
          conv2d_24_skip_comp <= 0;
          conv2d_24_skip_write_out <= 1;
          if(_maxi_read_req_idle) begin
            control_conv2d_24 <= control_conv2d_24_3;
          end 
        end
        control_conv2d_24_3: begin
          if(_maxi_read_idle) begin
            control_conv2d_24 <= control_conv2d_24_4;
          end 
        end
        control_conv2d_24_4: begin
          if(_maxi_read_req_idle) begin
            control_conv2d_24 <= control_conv2d_24_5;
          end 
        end
        control_conv2d_24_5: begin
          if(_maxi_read_idle) begin
            control_conv2d_24 <= control_conv2d_24_6;
          end 
        end
        control_conv2d_24_6: begin
          if(cparam_conv2d_24_data_stationary == 0) begin
            control_conv2d_24 <= control_conv2d_24_7;
          end 
          if(cparam_conv2d_24_data_stationary == 1) begin
            control_conv2d_24 <= control_conv2d_24_12;
          end 
        end
        control_conv2d_24_7: begin
          control_conv2d_24 <= control_conv2d_24_8;
          if(conv2d_24_skip_read_filter) begin
            control_conv2d_24 <= control_conv2d_24_11;
          end 
        end
        control_conv2d_24_8: begin
          if(_maxi_read_req_idle) begin
            control_conv2d_24 <= control_conv2d_24_9;
          end 
        end
        control_conv2d_24_9: begin
          if(_maxi_read_idle) begin
            control_conv2d_24 <= control_conv2d_24_10;
          end 
        end
        control_conv2d_24_10: begin
          control_conv2d_24 <= control_conv2d_24_11;
        end
        control_conv2d_24_11: begin
          if(cparam_conv2d_24_data_stationary == 0) begin
            control_conv2d_24 <= control_conv2d_24_12;
          end 
          if(cparam_conv2d_24_data_stationary == 1) begin
            control_conv2d_24 <= control_conv2d_24_24;
          end 
        end
        control_conv2d_24_12: begin
          control_conv2d_24 <= control_conv2d_24_13;
          if(conv2d_24_skip_read_act) begin
            control_conv2d_24 <= control_conv2d_24_23;
          end 
        end
        control_conv2d_24_13: begin
          control_conv2d_24 <= control_conv2d_24_14;
          if(conv2d_24_mux_dma_pad_mask_0 || !conv2d_24_mux_dma_flag_0) begin
            control_conv2d_24 <= control_conv2d_24_16;
          end 
        end
        control_conv2d_24_14: begin
          if(_maxi_read_req_idle) begin
            control_conv2d_24 <= control_conv2d_24_15;
          end 
        end
        control_conv2d_24_15: begin
          if(_maxi_read_idle) begin
            control_conv2d_24 <= control_conv2d_24_16;
          end 
        end
        control_conv2d_24_16: begin
          control_conv2d_24 <= control_conv2d_24_17;
          if(conv2d_24_mux_dma_pad_mask_1 || !conv2d_24_mux_dma_flag_1) begin
            control_conv2d_24 <= control_conv2d_24_19;
          end 
        end
        control_conv2d_24_17: begin
          if(_maxi_read_req_idle) begin
            control_conv2d_24 <= control_conv2d_24_18;
          end 
        end
        control_conv2d_24_18: begin
          if(_maxi_read_idle) begin
            control_conv2d_24 <= control_conv2d_24_19;
          end 
        end
        control_conv2d_24_19: begin
          control_conv2d_24 <= control_conv2d_24_20;
          if(conv2d_24_mux_dma_pad_mask_2 || !conv2d_24_mux_dma_flag_2) begin
            control_conv2d_24 <= control_conv2d_24_22;
          end 
        end
        control_conv2d_24_20: begin
          if(_maxi_read_req_idle) begin
            control_conv2d_24 <= control_conv2d_24_21;
          end 
        end
        control_conv2d_24_21: begin
          if(_maxi_read_idle) begin
            control_conv2d_24 <= control_conv2d_24_22;
          end 
        end
        control_conv2d_24_22: begin
          control_conv2d_24 <= control_conv2d_24_23;
        end
        control_conv2d_24_23: begin
          if(cparam_conv2d_24_data_stationary == 0) begin
            control_conv2d_24 <= control_conv2d_24_24;
          end 
          if(cparam_conv2d_24_data_stationary == 1) begin
            control_conv2d_24 <= control_conv2d_24_7;
          end 
        end
        control_conv2d_24_24: begin
          if(_maxi_write_idle) begin
            control_conv2d_24 <= control_conv2d_24_25;
          end 
        end
        control_conv2d_24_25: begin
          if(conv2d_24_comp_fsm == 0) begin
            control_conv2d_24 <= control_conv2d_24_26;
          end 
        end
        control_conv2d_24_26: begin
          control_conv2d_24 <= control_conv2d_24_27;
          if(conv2d_24_skip_write_out) begin
            control_conv2d_24 <= control_conv2d_24_32;
          end 
          if((cparam_conv2d_24_data_stationary == 1) && (conv2d_24_prev_och_count < cparam_conv2d_24_max_och_count)) begin
            control_conv2d_24 <= control_conv2d_24_32;
          end 
        end
        control_conv2d_24_27: begin
          if(conv2d_24_sync_comp_count >= conv2d_24_sync_out_count + cparam_conv2d_24_inc_sync_out) begin
            control_conv2d_24 <= control_conv2d_24_28;
          end 
        end
        control_conv2d_24_28: begin
          if(!conv2d_24_dma_out_mask_0) begin
            control_conv2d_24 <= control_conv2d_24_29;
          end 
          if(conv2d_24_dma_out_mask_0) begin
            control_conv2d_24 <= control_conv2d_24_30;
          end 
        end
        control_conv2d_24_29: begin
          if(_maxi_write_req_idle) begin
            control_conv2d_24 <= control_conv2d_24_30;
          end 
        end
        control_conv2d_24_30: begin
          control_conv2d_24 <= control_conv2d_24_31;
        end
        control_conv2d_24_31: begin
          conv2d_24_write_count <= conv2d_24_write_count + 1;
          if(conv2d_24_out_ram_select == 0) begin
            conv2d_24_out_laddr_offset <= conv2d_24_out_laddr_offset + conv2d_24_next_out_write_size;
          end 
          if((cparam_conv2d_24_data_stationary == 0) && !cparam_conv2d_24_keep_filter) begin
            conv2d_24_out_base_offset_col <= conv2d_24_out_base_offset_col + cparam_conv2d_24_out_col_step;
            conv2d_24_out_col_count <= conv2d_24_out_col_count + 1;
          end 
          conv2d_24_out_ram_select <= conv2d_24_out_ram_select + 1;
          if(conv2d_24_out_ram_select == 0) begin
            conv2d_24_out_ram_select <= 0;
          end 
          conv2d_24_sync_out_count <= conv2d_24_sync_out_count + cparam_conv2d_24_inc_sync_out;
          if((cparam_conv2d_24_data_stationary == 0) && !cparam_conv2d_24_keep_filter && (conv2d_24_write_count >= cparam_conv2d_24_out_num_col - 1) || (cparam_conv2d_24_data_stationary == 0) && cparam_conv2d_24_keep_filter || (cparam_conv2d_24_data_stationary == 1)) begin
            conv2d_24_sync_out_count <= conv2d_24_sync_out_count + (cparam_conv2d_24_inc_sync_out + cparam_conv2d_24_inc_sync_out_res);
          end 
          if((cparam_conv2d_24_data_stationary == 0) && !cparam_conv2d_24_keep_filter) begin
            control_conv2d_24 <= control_conv2d_24_26;
          end 
          if((cparam_conv2d_24_data_stationary == 0) && !cparam_conv2d_24_keep_filter && (conv2d_24_write_count >= cparam_conv2d_24_out_num_col - 1) || (cparam_conv2d_24_data_stationary == 0) && cparam_conv2d_24_keep_filter || (cparam_conv2d_24_data_stationary == 1)) begin
            control_conv2d_24 <= control_conv2d_24_32;
          end 
        end
        control_conv2d_24_32: begin
          if(conv2d_24_update_filter) begin
            conv2d_24_filter_base_offset <= conv2d_24_filter_base_offset + cparam_conv2d_24_filter_base_step;
          end 
          if((cparam_conv2d_24_data_stationary == 1) && (conv2d_24_och_count >= cparam_conv2d_24_max_och_count)) begin
            conv2d_24_filter_base_offset <= 0;
          end 
          if(conv2d_24_update_filter) begin
            conv2d_24_och_count <= conv2d_24_och_count + cparam_conv2d_24_och_count_step;
          end 
          if((cparam_conv2d_24_data_stationary == 1) && (conv2d_24_och_count >= cparam_conv2d_24_max_och_count)) begin
            conv2d_24_och_count <= 0;
          end 
          if(conv2d_24_update_filter) begin
            conv2d_24_filter_page_comp_offset <= conv2d_24_filter_page_comp_offset + cparam_conv2d_24_filter_read_step;
            conv2d_24_filter_page_dma_offset <= conv2d_24_filter_page_dma_offset + cparam_conv2d_24_filter_read_step;
          end 
          if(conv2d_24_update_filter && (conv2d_24_filter_page_comp_offset + cparam_conv2d_24_filter_read_step + cparam_conv2d_24_filter_read_step > 4096)) begin
            conv2d_24_filter_page_comp_offset <= 0;
            conv2d_24_filter_page_dma_offset <= 0;
          end 
          if(conv2d_24_update_act) begin
            conv2d_24_act_base_offset_row <= conv2d_24_act_base_offset_row + cparam_conv2d_24_act_row_step;
          end 
          if(conv2d_24_update_act && (conv2d_24_row_count >= cparam_conv2d_24_max_row_count)) begin
            conv2d_24_act_base_offset_row <= 0;
            conv2d_24_act_base_offset_bat <= conv2d_24_act_base_offset_bat + cparam_conv2d_24_act_bat_step;
          end 
          if(conv2d_24_update_act && (conv2d_24_row_count >= cparam_conv2d_24_max_row_count) && (conv2d_24_bat_count >= cparam_conv2d_24_max_bat_count)) begin
            conv2d_24_act_base_offset_bat <= 0;
          end 
          if(!conv2d_24_update_act) begin
            conv2d_24_dma_flag_0 <= 0;
          end 
          if(conv2d_24_update_act) begin
            conv2d_24_dma_flag_0 <= cparam_conv2d_24_dma_flag_conds_0;
          end 
          if(conv2d_24_update_act && (conv2d_24_row_count >= cparam_conv2d_24_max_row_count)) begin
            conv2d_24_dma_flag_0 <= 1;
          end 
          if(!conv2d_24_update_act) begin
            conv2d_24_dma_flag_1 <= 0;
          end 
          if(conv2d_24_update_act) begin
            conv2d_24_dma_flag_1 <= cparam_conv2d_24_dma_flag_conds_1;
          end 
          if(conv2d_24_update_act && (conv2d_24_row_count >= cparam_conv2d_24_max_row_count)) begin
            conv2d_24_dma_flag_1 <= 1;
          end 
          if(!conv2d_24_update_act) begin
            conv2d_24_dma_flag_2 <= 0;
          end 
          if(conv2d_24_update_act) begin
            conv2d_24_dma_flag_2 <= cparam_conv2d_24_dma_flag_conds_2;
          end 
          if(conv2d_24_update_act && (conv2d_24_row_count >= cparam_conv2d_24_max_row_count)) begin
            conv2d_24_dma_flag_2 <= 1;
          end 
          if(conv2d_24_update_act) begin
            conv2d_24_row_count <= conv2d_24_row_count + cparam_conv2d_24_stride_row_par_row;
          end 
          if(conv2d_24_update_act && (conv2d_24_row_count >= cparam_conv2d_24_max_row_count)) begin
            conv2d_24_row_count <= 0;
            conv2d_24_bat_count <= conv2d_24_bat_count + 1;
          end 
          if(conv2d_24_update_act && (conv2d_24_row_count >= cparam_conv2d_24_max_row_count) && (conv2d_24_bat_count >= cparam_conv2d_24_max_bat_count)) begin
            conv2d_24_bat_count <= 0;
          end 
          if(conv2d_24_update_act && (cparam_conv2d_24_stride_row_par_row < 3)) begin
            conv2d_24_row_select <= conv2d_24_row_select + cparam_conv2d_24_stride_row_par_row;
            conv2d_24_prev_row_select <= conv2d_24_row_select;
          end 
          if(conv2d_24_update_act && (cparam_conv2d_24_stride_row_par_row < 3) && (conv2d_24_row_select + cparam_conv2d_24_stride_row_par_row >= 3)) begin
            conv2d_24_row_select <= conv2d_24_row_select - (3 - cparam_conv2d_24_stride_row_par_row);
            conv2d_24_prev_row_select <= conv2d_24_row_select;
          end 
          if(conv2d_24_update_act && !(cparam_conv2d_24_stride_row_par_row < 3)) begin
            conv2d_24_row_select <= 0;
            conv2d_24_prev_row_select <= 0;
          end 
          if(conv2d_24_update_act && (conv2d_24_row_count >= cparam_conv2d_24_max_row_count)) begin
            conv2d_24_row_select <= 0;
            conv2d_24_prev_row_select <= 0;
          end 
          if(conv2d_24_update_act && conv2d_24_mux_next_dma_flag_0) begin
            conv2d_24_act_page_comp_offset_0 <= conv2d_24_act_page_comp_offset_0 + cparam_conv2d_24_act_read_step;
            conv2d_24_act_page_dma_offset_0 <= conv2d_24_act_page_dma_offset_0 + cparam_conv2d_24_act_read_step;
          end 
          if(conv2d_24_update_act && conv2d_24_mux_next_dma_flag_0 && (conv2d_24_act_page_comp_offset_0 + cparam_conv2d_24_act_read_step + cparam_conv2d_24_act_read_step > 16384)) begin
            conv2d_24_act_page_comp_offset_0 <= 0;
            conv2d_24_act_page_dma_offset_0 <= 0;
          end 
          if((cparam_conv2d_24_data_stationary == 0) && (conv2d_24_row_count >= cparam_conv2d_24_max_row_count) && (conv2d_24_bat_count >= cparam_conv2d_24_max_bat_count) && cparam_conv2d_24_keep_input) begin
            conv2d_24_act_page_comp_offset_0 <= 0;
            conv2d_24_act_page_dma_offset_0 <= 0;
          end 
          if(conv2d_24_update_act && conv2d_24_mux_next_dma_flag_1) begin
            conv2d_24_act_page_comp_offset_1 <= conv2d_24_act_page_comp_offset_1 + cparam_conv2d_24_act_read_step;
            conv2d_24_act_page_dma_offset_1 <= conv2d_24_act_page_dma_offset_1 + cparam_conv2d_24_act_read_step;
          end 
          if(conv2d_24_update_act && conv2d_24_mux_next_dma_flag_1 && (conv2d_24_act_page_comp_offset_1 + cparam_conv2d_24_act_read_step + cparam_conv2d_24_act_read_step > 16384)) begin
            conv2d_24_act_page_comp_offset_1 <= 0;
            conv2d_24_act_page_dma_offset_1 <= 0;
          end 
          if((cparam_conv2d_24_data_stationary == 0) && (conv2d_24_row_count >= cparam_conv2d_24_max_row_count) && (conv2d_24_bat_count >= cparam_conv2d_24_max_bat_count) && cparam_conv2d_24_keep_input) begin
            conv2d_24_act_page_comp_offset_1 <= 0;
            conv2d_24_act_page_dma_offset_1 <= 0;
          end 
          if(conv2d_24_update_act && conv2d_24_mux_next_dma_flag_2) begin
            conv2d_24_act_page_comp_offset_2 <= conv2d_24_act_page_comp_offset_2 + cparam_conv2d_24_act_read_step;
            conv2d_24_act_page_dma_offset_2 <= conv2d_24_act_page_dma_offset_2 + cparam_conv2d_24_act_read_step;
          end 
          if(conv2d_24_update_act && conv2d_24_mux_next_dma_flag_2 && (conv2d_24_act_page_comp_offset_2 + cparam_conv2d_24_act_read_step + cparam_conv2d_24_act_read_step > 16384)) begin
            conv2d_24_act_page_comp_offset_2 <= 0;
            conv2d_24_act_page_dma_offset_2 <= 0;
          end 
          if((cparam_conv2d_24_data_stationary == 0) && (conv2d_24_row_count >= cparam_conv2d_24_max_row_count) && (conv2d_24_bat_count >= cparam_conv2d_24_max_bat_count) && cparam_conv2d_24_keep_input) begin
            conv2d_24_act_page_comp_offset_2 <= 0;
            conv2d_24_act_page_dma_offset_2 <= 0;
          end 
          conv2d_24_next_out_write_size <= (conv2d_24_och_count >= cparam_conv2d_24_max_och_count)? cparam_conv2d_24_out_write_size_res : cparam_conv2d_24_out_write_size;
          if(!conv2d_24_skip_write_out) begin
            conv2d_24_write_count <= 0;
            conv2d_24_out_laddr_offset <= 0;
            conv2d_24_out_ram_select <= 0;
          end 
          if((cparam_conv2d_24_data_stationary == 0) && !conv2d_24_skip_write_out) begin
            conv2d_24_out_base_offset_col <= 0;
            conv2d_24_out_base_offset_row <= conv2d_24_out_base_offset_row + cparam_conv2d_24_out_row_step;
            conv2d_24_out_col_count <= 0;
            conv2d_24_out_row_count <= conv2d_24_out_row_count + 1;
          end 
          if((cparam_conv2d_24_data_stationary == 0) && !conv2d_24_skip_write_out && (conv2d_24_prev_row_count >= cparam_conv2d_24_max_row_count)) begin
            conv2d_24_out_base_offset_row <= 0;
            conv2d_24_out_base_offset_bat <= conv2d_24_out_base_offset_bat + cparam_conv2d_24_out_bat_step;
            conv2d_24_out_row_count <= 0;
          end 
          if((cparam_conv2d_24_data_stationary == 0) && !conv2d_24_skip_write_out && (conv2d_24_prev_row_count >= cparam_conv2d_24_max_row_count) && (conv2d_24_prev_bat_count >= cparam_conv2d_24_max_bat_count)) begin
            conv2d_24_out_base_offset_bat <= 0;
            conv2d_24_out_base_offset_och <= conv2d_24_out_base_offset_och + cparam_conv2d_24_out_och_step;
          end 
          if((cparam_conv2d_24_data_stationary == 1) && (conv2d_24_prev_och_count >= cparam_conv2d_24_max_och_count) && !conv2d_24_skip_write_out) begin
            conv2d_24_out_base_offset_row <= conv2d_24_out_base_offset_row + cparam_conv2d_24_out_row_step;
          end 
          if((cparam_conv2d_24_data_stationary == 0) && !conv2d_24_out_page) begin
            conv2d_24_out_page_comp_offset <= 1024;
            conv2d_24_out_page_dma_offset <= 0;
            conv2d_24_out_page <= 1;
          end 
          if((cparam_conv2d_24_data_stationary == 0) && conv2d_24_out_page) begin
            conv2d_24_out_page_comp_offset <= 0;
            conv2d_24_out_page_dma_offset <= 1024;
            conv2d_24_out_page <= 0;
          end 
          if((cparam_conv2d_24_data_stationary == 1) && (conv2d_24_och_count >= cparam_conv2d_24_max_och_count) && !conv2d_24_out_page) begin
            conv2d_24_out_page_comp_offset <= 1024;
            conv2d_24_out_page_dma_offset <= 0;
            conv2d_24_out_page <= 1;
          end 
          if((cparam_conv2d_24_data_stationary == 1) && (conv2d_24_och_count >= cparam_conv2d_24_max_och_count) && conv2d_24_out_page) begin
            conv2d_24_out_page_comp_offset <= 0;
            conv2d_24_out_page_dma_offset <= 1024;
            conv2d_24_out_page <= 0;
          end 
          conv2d_24_prev_row_count <= conv2d_24_row_count;
          conv2d_24_prev_bat_count <= conv2d_24_bat_count;
          conv2d_24_prev_och_count <= conv2d_24_och_count;
          if((conv2d_24_row_count >= cparam_conv2d_24_max_row_count) && (conv2d_24_bat_count >= cparam_conv2d_24_max_bat_count) && (conv2d_24_och_count >= cparam_conv2d_24_max_och_count)) begin
            conv2d_24_skip_read_filter <= 1;
          end 
          if((cparam_conv2d_24_data_stationary == 1) && cparam_conv2d_24_keep_filter) begin
            conv2d_24_skip_read_filter <= 1;
          end 
          if((conv2d_24_row_count >= cparam_conv2d_24_max_row_count) && (conv2d_24_bat_count >= cparam_conv2d_24_max_bat_count) && (conv2d_24_och_count >= cparam_conv2d_24_max_och_count)) begin
            conv2d_24_skip_read_act <= 1;
          end 
          if((cparam_conv2d_24_data_stationary == 0) && (conv2d_24_row_count >= cparam_conv2d_24_max_row_count) && (conv2d_24_bat_count >= cparam_conv2d_24_max_bat_count) && cparam_conv2d_24_keep_input) begin
            conv2d_24_skip_read_act <= 1;
          end 
          if((conv2d_24_row_count >= cparam_conv2d_24_max_row_count) && (conv2d_24_bat_count >= cparam_conv2d_24_max_bat_count) && (conv2d_24_och_count >= cparam_conv2d_24_max_och_count)) begin
            conv2d_24_skip_comp <= 1;
          end 
          if(conv2d_24_skip_write_out && (conv2d_24_prev_row_count == 0) && (conv2d_24_prev_bat_count == 0) && (conv2d_24_prev_och_count == 0)) begin
            conv2d_24_skip_write_out <= 0;
          end 
          if(cparam_conv2d_24_data_stationary == 0) begin
            control_conv2d_24 <= control_conv2d_24_12;
          end 
          if((cparam_conv2d_24_data_stationary == 0) && (conv2d_24_row_count >= cparam_conv2d_24_max_row_count) && (conv2d_24_bat_count >= cparam_conv2d_24_max_bat_count)) begin
            control_conv2d_24 <= control_conv2d_24_7;
          end 
          if(cparam_conv2d_24_data_stationary == 1) begin
            control_conv2d_24 <= control_conv2d_24_7;
          end 
          if((cparam_conv2d_24_data_stationary == 1) && (conv2d_24_och_count >= cparam_conv2d_24_max_och_count)) begin
            control_conv2d_24 <= control_conv2d_24_12;
          end 
          if(!conv2d_24_skip_write_out && (conv2d_24_prev_och_count >= cparam_conv2d_24_max_och_count) && (conv2d_24_prev_row_count >= cparam_conv2d_24_max_row_count) && (conv2d_24_prev_bat_count >= cparam_conv2d_24_max_bat_count)) begin
            control_conv2d_24 <= control_conv2d_24_33;
          end 
        end
        control_conv2d_24_33: begin
          if(_maxi_write_idle && !_maxi_has_outstanding_write) begin
            control_conv2d_24 <= control_conv2d_24_34;
          end 
        end
        control_conv2d_24_34: begin
          if(main_fsm == 14) begin
            _control_conv2d_24_called <= 0;
          end 
          if(main_fsm == 31) begin
            _control_conv2d_24_called <= 0;
          end 
          if(main_fsm == 48) begin
            _control_conv2d_24_called <= 0;
          end 
          if(main_fsm == 58) begin
            _control_conv2d_24_called <= 0;
          end 
          if(main_fsm == 75) begin
            _control_conv2d_24_called <= 0;
          end 
          if(main_fsm == 85) begin
            _control_conv2d_24_called <= 0;
          end 
          if(main_fsm == 102) begin
            _control_conv2d_24_called <= 0;
          end 
          if(main_fsm == 112) begin
            _control_conv2d_24_called <= 0;
          end 
          if(main_fsm == 14) begin
            control_conv2d_24 <= control_conv2d_24_init;
          end 
          if(main_fsm == 31) begin
            control_conv2d_24 <= control_conv2d_24_init;
          end 
          if(main_fsm == 48) begin
            control_conv2d_24 <= control_conv2d_24_init;
          end 
          if(main_fsm == 58) begin
            control_conv2d_24 <= control_conv2d_24_init;
          end 
          if(main_fsm == 75) begin
            control_conv2d_24 <= control_conv2d_24_init;
          end 
          if(main_fsm == 85) begin
            control_conv2d_24 <= control_conv2d_24_init;
          end 
          if(main_fsm == 102) begin
            control_conv2d_24 <= control_conv2d_24_init;
          end 
          if(main_fsm == 112) begin
            control_conv2d_24 <= control_conv2d_24_init;
          end 
        end
      endcase
    end
  end

  localparam _maxi_read_req_fsm_1 = 1;

  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      _maxi_read_req_fsm <= _maxi_read_req_fsm_init;
      _maxi_read_cont <= 0;
    end else begin
      case(_maxi_read_req_fsm)
        _maxi_read_req_fsm_init: begin
          if((_maxi_read_req_fsm == 0) && (_maxi_read_start || _maxi_read_cont) && !_maxi_read_req_fifo_almost_full) begin
            _maxi_read_req_fsm <= _maxi_read_req_fsm_1;
          end 
        end
        _maxi_read_req_fsm_1: begin
          if(maxi_arready || !maxi_arvalid) begin
            _maxi_read_cont <= 1;
          end 
          if((maxi_arready || !maxi_arvalid) && (_maxi_read_global_size == 0)) begin
            _maxi_read_cont <= 0;
          end 
          if(maxi_arready || !maxi_arvalid) begin
            _maxi_read_req_fsm <= _maxi_read_req_fsm_init;
          end 
        end
      endcase
    end
  end

  localparam _maxi_read_data_fsm_1 = 1;
  localparam _maxi_read_data_fsm_2 = 2;

  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
    end else begin
      case(_maxi_read_data_fsm)
        _maxi_read_data_fsm_init: begin
          if(!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
          if(!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 2)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
          if(!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 3)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
          if(!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 4)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
          if(!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 5)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
          if(!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 6)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
          if(!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 7)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
          if(!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 8)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
          if(!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 9)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
        end
        _maxi_read_data_fsm_1: begin
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
        end
        _maxi_read_data_fsm_2: begin
          if(_maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
          if(_maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
          if(_maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
          if(_maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
          if(_maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
          if(_maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
          if(_maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
          if(_maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
          if(_maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_0_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_0 <= write_burst_fsm_0_init;
      write_burst_addr_76 <= 0;
      write_burst_stride_77 <= 0;
      write_burst_length_78 <= 0;
      write_burst_done_79 <= 0;
    end else begin
      case(write_burst_fsm_0)
        write_burst_fsm_0_init: begin
          write_burst_addr_76 <= _maxi_read_local_addr_buf;
          write_burst_stride_77 <= _maxi_read_local_stride_buf;
          write_burst_length_78 <= _maxi_read_local_size_buf;
          write_burst_done_79 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 1) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_fsm_0 <= write_burst_fsm_0_1;
          end 
        end
        write_burst_fsm_0_1: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_addr_76 <= write_burst_addr_76 + write_burst_stride_77;
            write_burst_length_78 <= write_burst_length_78 - 1;
            write_burst_done_79 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_length_78 <= 1)) begin
            write_burst_done_79 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_done_79 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_length_78 <= 1)) begin
            write_burst_fsm_0 <= write_burst_fsm_0_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_fsm_0 <= write_burst_fsm_0_init;
          end 
          if(0) begin
            write_burst_fsm_0 <= write_burst_fsm_0_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_1_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_1 <= write_burst_packed_fsm_1_init;
      write_burst_packed_addr_85 <= 0;
      write_burst_packed_stride_86 <= 0;
      write_burst_packed_length_87 <= 0;
      write_burst_packed_done_88 <= 0;
    end else begin
      case(write_burst_packed_fsm_1)
        write_burst_packed_fsm_1_init: begin
          write_burst_packed_addr_85 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_86 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_87 <= _maxi_read_local_size_buf;
          write_burst_packed_done_88 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 2) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_1 <= write_burst_packed_fsm_1_1;
          end 
        end
        write_burst_packed_fsm_1_1: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_packed_addr_85 <= write_burst_packed_addr_85 + write_burst_packed_stride_86;
            write_burst_packed_length_87 <= write_burst_packed_length_87 - 1;
            write_burst_packed_done_88 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_packed_length_87 <= 1)) begin
            write_burst_packed_done_88 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_packed_done_88 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_packed_length_87 <= 1)) begin
            write_burst_packed_fsm_1 <= write_burst_packed_fsm_1_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_packed_fsm_1 <= write_burst_packed_fsm_1_init;
          end 
          if(0) begin
            write_burst_packed_fsm_1 <= write_burst_packed_fsm_1_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_2_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_2 <= write_burst_packed_fsm_2_init;
      write_burst_packed_addr_107 <= 0;
      write_burst_packed_stride_108 <= 0;
      write_burst_packed_length_109 <= 0;
      write_burst_packed_done_110 <= 0;
    end else begin
      case(write_burst_packed_fsm_2)
        write_burst_packed_fsm_2_init: begin
          write_burst_packed_addr_107 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_108 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_109 <= _maxi_read_local_size_buf;
          write_burst_packed_done_110 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_2 <= write_burst_packed_fsm_2_1;
          end 
        end
        write_burst_packed_fsm_2_1: begin
          if(write_burst_block_ram_wvalid_105) begin
            write_burst_packed_addr_107 <= write_burst_packed_addr_107 + write_burst_packed_stride_108;
            write_burst_packed_length_109 <= write_burst_packed_length_109 - 1;
            write_burst_packed_done_110 <= 0;
          end 
          if(write_burst_block_ram_wvalid_105 && (write_burst_packed_length_109 <= 1)) begin
            write_burst_packed_done_110 <= 1;
          end 
          if(write_burst_block_ram_wvalid_105 && 0) begin
            write_burst_packed_done_110 <= 1;
          end 
          if(write_burst_block_ram_wvalid_105 && (write_burst_packed_length_109 <= 1)) begin
            write_burst_packed_fsm_2 <= write_burst_packed_fsm_2_init;
          end 
          if(write_burst_block_ram_wvalid_105 && 0) begin
            write_burst_packed_fsm_2 <= write_burst_packed_fsm_2_init;
          end 
          if(write_burst_block_ram_wquit_106) begin
            write_burst_packed_fsm_2 <= write_burst_packed_fsm_2_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_3_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_3 <= write_burst_packed_fsm_3_init;
      write_burst_packed_addr_121 <= 0;
      write_burst_packed_stride_122 <= 0;
      write_burst_packed_length_123 <= 0;
      write_burst_packed_done_124 <= 0;
    end else begin
      case(write_burst_packed_fsm_3)
        write_burst_packed_fsm_3_init: begin
          write_burst_packed_addr_121 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_122 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_123 <= _maxi_read_local_size_buf;
          write_burst_packed_done_124 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_3 <= write_burst_packed_fsm_3_1;
          end 
        end
        write_burst_packed_fsm_3_1: begin
          if(write_burst_block_ram_wvalid_119) begin
            write_burst_packed_addr_121 <= write_burst_packed_addr_121 + write_burst_packed_stride_122;
            write_burst_packed_length_123 <= write_burst_packed_length_123 - 1;
            write_burst_packed_done_124 <= 0;
          end 
          if(write_burst_block_ram_wvalid_119 && (write_burst_packed_length_123 <= 1)) begin
            write_burst_packed_done_124 <= 1;
          end 
          if(write_burst_block_ram_wvalid_119 && 0) begin
            write_burst_packed_done_124 <= 1;
          end 
          if(write_burst_block_ram_wvalid_119 && (write_burst_packed_length_123 <= 1)) begin
            write_burst_packed_fsm_3 <= write_burst_packed_fsm_3_init;
          end 
          if(write_burst_block_ram_wvalid_119 && 0) begin
            write_burst_packed_fsm_3 <= write_burst_packed_fsm_3_init;
          end 
          if(write_burst_block_ram_wquit_120) begin
            write_burst_packed_fsm_3 <= write_burst_packed_fsm_3_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_4_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_4 <= write_burst_packed_fsm_4_init;
      write_burst_packed_addr_135 <= 0;
      write_burst_packed_stride_136 <= 0;
      write_burst_packed_length_137 <= 0;
      write_burst_packed_done_138 <= 0;
    end else begin
      case(write_burst_packed_fsm_4)
        write_burst_packed_fsm_4_init: begin
          write_burst_packed_addr_135 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_136 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_137 <= _maxi_read_local_size_buf;
          write_burst_packed_done_138 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_4 <= write_burst_packed_fsm_4_1;
          end 
        end
        write_burst_packed_fsm_4_1: begin
          if(write_burst_block_ram_wvalid_133) begin
            write_burst_packed_addr_135 <= write_burst_packed_addr_135 + write_burst_packed_stride_136;
            write_burst_packed_length_137 <= write_burst_packed_length_137 - 1;
            write_burst_packed_done_138 <= 0;
          end 
          if(write_burst_block_ram_wvalid_133 && (write_burst_packed_length_137 <= 1)) begin
            write_burst_packed_done_138 <= 1;
          end 
          if(write_burst_block_ram_wvalid_133 && 0) begin
            write_burst_packed_done_138 <= 1;
          end 
          if(write_burst_block_ram_wvalid_133 && (write_burst_packed_length_137 <= 1)) begin
            write_burst_packed_fsm_4 <= write_burst_packed_fsm_4_init;
          end 
          if(write_burst_block_ram_wvalid_133 && 0) begin
            write_burst_packed_fsm_4 <= write_burst_packed_fsm_4_init;
          end 
          if(write_burst_block_ram_wquit_134) begin
            write_burst_packed_fsm_4 <= write_burst_packed_fsm_4_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_5_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_5 <= write_burst_packed_fsm_5_init;
      write_burst_packed_addr_149 <= 0;
      write_burst_packed_stride_150 <= 0;
      write_burst_packed_length_151 <= 0;
      write_burst_packed_done_152 <= 0;
    end else begin
      case(write_burst_packed_fsm_5)
        write_burst_packed_fsm_5_init: begin
          write_burst_packed_addr_149 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_150 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_151 <= _maxi_read_local_size_buf;
          write_burst_packed_done_152 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_5 <= write_burst_packed_fsm_5_1;
          end 
        end
        write_burst_packed_fsm_5_1: begin
          if(write_burst_block_ram_wvalid_147) begin
            write_burst_packed_addr_149 <= write_burst_packed_addr_149 + write_burst_packed_stride_150;
            write_burst_packed_length_151 <= write_burst_packed_length_151 - 1;
            write_burst_packed_done_152 <= 0;
          end 
          if(write_burst_block_ram_wvalid_147 && (write_burst_packed_length_151 <= 1)) begin
            write_burst_packed_done_152 <= 1;
          end 
          if(write_burst_block_ram_wvalid_147 && 0) begin
            write_burst_packed_done_152 <= 1;
          end 
          if(write_burst_block_ram_wvalid_147 && (write_burst_packed_length_151 <= 1)) begin
            write_burst_packed_fsm_5 <= write_burst_packed_fsm_5_init;
          end 
          if(write_burst_block_ram_wvalid_147 && 0) begin
            write_burst_packed_fsm_5 <= write_burst_packed_fsm_5_init;
          end 
          if(write_burst_block_ram_wquit_148) begin
            write_burst_packed_fsm_5 <= write_burst_packed_fsm_5_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_6_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_6 <= write_burst_packed_fsm_6_init;
      write_burst_packed_addr_163 <= 0;
      write_burst_packed_stride_164 <= 0;
      write_burst_packed_length_165 <= 0;
      write_burst_packed_done_166 <= 0;
    end else begin
      case(write_burst_packed_fsm_6)
        write_burst_packed_fsm_6_init: begin
          write_burst_packed_addr_163 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_164 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_165 <= _maxi_read_local_size_buf;
          write_burst_packed_done_166 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_6 <= write_burst_packed_fsm_6_1;
          end 
        end
        write_burst_packed_fsm_6_1: begin
          if(write_burst_block_ram_wvalid_161) begin
            write_burst_packed_addr_163 <= write_burst_packed_addr_163 + write_burst_packed_stride_164;
            write_burst_packed_length_165 <= write_burst_packed_length_165 - 1;
            write_burst_packed_done_166 <= 0;
          end 
          if(write_burst_block_ram_wvalid_161 && (write_burst_packed_length_165 <= 1)) begin
            write_burst_packed_done_166 <= 1;
          end 
          if(write_burst_block_ram_wvalid_161 && 0) begin
            write_burst_packed_done_166 <= 1;
          end 
          if(write_burst_block_ram_wvalid_161 && (write_burst_packed_length_165 <= 1)) begin
            write_burst_packed_fsm_6 <= write_burst_packed_fsm_6_init;
          end 
          if(write_burst_block_ram_wvalid_161 && 0) begin
            write_burst_packed_fsm_6 <= write_burst_packed_fsm_6_init;
          end 
          if(write_burst_block_ram_wquit_162) begin
            write_burst_packed_fsm_6 <= write_burst_packed_fsm_6_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_7_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_7 <= write_burst_packed_fsm_7_init;
      write_burst_packed_addr_177 <= 0;
      write_burst_packed_stride_178 <= 0;
      write_burst_packed_length_179 <= 0;
      write_burst_packed_done_180 <= 0;
    end else begin
      case(write_burst_packed_fsm_7)
        write_burst_packed_fsm_7_init: begin
          write_burst_packed_addr_177 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_178 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_179 <= _maxi_read_local_size_buf;
          write_burst_packed_done_180 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_7 <= write_burst_packed_fsm_7_1;
          end 
        end
        write_burst_packed_fsm_7_1: begin
          if(write_burst_block_ram_wvalid_175) begin
            write_burst_packed_addr_177 <= write_burst_packed_addr_177 + write_burst_packed_stride_178;
            write_burst_packed_length_179 <= write_burst_packed_length_179 - 1;
            write_burst_packed_done_180 <= 0;
          end 
          if(write_burst_block_ram_wvalid_175 && (write_burst_packed_length_179 <= 1)) begin
            write_burst_packed_done_180 <= 1;
          end 
          if(write_burst_block_ram_wvalid_175 && 0) begin
            write_burst_packed_done_180 <= 1;
          end 
          if(write_burst_block_ram_wvalid_175 && (write_burst_packed_length_179 <= 1)) begin
            write_burst_packed_fsm_7 <= write_burst_packed_fsm_7_init;
          end 
          if(write_burst_block_ram_wvalid_175 && 0) begin
            write_burst_packed_fsm_7 <= write_burst_packed_fsm_7_init;
          end 
          if(write_burst_block_ram_wquit_176) begin
            write_burst_packed_fsm_7 <= write_burst_packed_fsm_7_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_8_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_8 <= write_burst_packed_fsm_8_init;
      write_burst_packed_addr_191 <= 0;
      write_burst_packed_stride_192 <= 0;
      write_burst_packed_length_193 <= 0;
      write_burst_packed_done_194 <= 0;
    end else begin
      case(write_burst_packed_fsm_8)
        write_burst_packed_fsm_8_init: begin
          write_burst_packed_addr_191 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_192 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_193 <= _maxi_read_local_size_buf;
          write_burst_packed_done_194 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_8 <= write_burst_packed_fsm_8_1;
          end 
        end
        write_burst_packed_fsm_8_1: begin
          if(write_burst_block_ram_wvalid_189) begin
            write_burst_packed_addr_191 <= write_burst_packed_addr_191 + write_burst_packed_stride_192;
            write_burst_packed_length_193 <= write_burst_packed_length_193 - 1;
            write_burst_packed_done_194 <= 0;
          end 
          if(write_burst_block_ram_wvalid_189 && (write_burst_packed_length_193 <= 1)) begin
            write_burst_packed_done_194 <= 1;
          end 
          if(write_burst_block_ram_wvalid_189 && 0) begin
            write_burst_packed_done_194 <= 1;
          end 
          if(write_burst_block_ram_wvalid_189 && (write_burst_packed_length_193 <= 1)) begin
            write_burst_packed_fsm_8 <= write_burst_packed_fsm_8_init;
          end 
          if(write_burst_block_ram_wvalid_189 && 0) begin
            write_burst_packed_fsm_8 <= write_burst_packed_fsm_8_init;
          end 
          if(write_burst_block_ram_wquit_190) begin
            write_burst_packed_fsm_8 <= write_burst_packed_fsm_8_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_9_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_9 <= write_burst_packed_fsm_9_init;
      write_burst_packed_addr_205 <= 0;
      write_burst_packed_stride_206 <= 0;
      write_burst_packed_length_207 <= 0;
      write_burst_packed_done_208 <= 0;
    end else begin
      case(write_burst_packed_fsm_9)
        write_burst_packed_fsm_9_init: begin
          write_burst_packed_addr_205 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_206 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_207 <= _maxi_read_local_size_buf;
          write_burst_packed_done_208 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_9 <= write_burst_packed_fsm_9_1;
          end 
        end
        write_burst_packed_fsm_9_1: begin
          if(write_burst_block_ram_wvalid_203) begin
            write_burst_packed_addr_205 <= write_burst_packed_addr_205 + write_burst_packed_stride_206;
            write_burst_packed_length_207 <= write_burst_packed_length_207 - 1;
            write_burst_packed_done_208 <= 0;
          end 
          if(write_burst_block_ram_wvalid_203 && (write_burst_packed_length_207 <= 1)) begin
            write_burst_packed_done_208 <= 1;
          end 
          if(write_burst_block_ram_wvalid_203 && 0) begin
            write_burst_packed_done_208 <= 1;
          end 
          if(write_burst_block_ram_wvalid_203 && (write_burst_packed_length_207 <= 1)) begin
            write_burst_packed_fsm_9 <= write_burst_packed_fsm_9_init;
          end 
          if(write_burst_block_ram_wvalid_203 && 0) begin
            write_burst_packed_fsm_9 <= write_burst_packed_fsm_9_init;
          end 
          if(write_burst_block_ram_wquit_204) begin
            write_burst_packed_fsm_9 <= write_burst_packed_fsm_9_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_10_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_10 <= write_burst_packed_fsm_10_init;
      write_burst_packed_addr_219 <= 0;
      write_burst_packed_stride_220 <= 0;
      write_burst_packed_length_221 <= 0;
      write_burst_packed_done_222 <= 0;
    end else begin
      case(write_burst_packed_fsm_10)
        write_burst_packed_fsm_10_init: begin
          write_burst_packed_addr_219 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_220 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_221 <= _maxi_read_local_size_buf;
          write_burst_packed_done_222 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_10 <= write_burst_packed_fsm_10_1;
          end 
        end
        write_burst_packed_fsm_10_1: begin
          if(write_burst_block_ram_wvalid_217) begin
            write_burst_packed_addr_219 <= write_burst_packed_addr_219 + write_burst_packed_stride_220;
            write_burst_packed_length_221 <= write_burst_packed_length_221 - 1;
            write_burst_packed_done_222 <= 0;
          end 
          if(write_burst_block_ram_wvalid_217 && (write_burst_packed_length_221 <= 1)) begin
            write_burst_packed_done_222 <= 1;
          end 
          if(write_burst_block_ram_wvalid_217 && 0) begin
            write_burst_packed_done_222 <= 1;
          end 
          if(write_burst_block_ram_wvalid_217 && (write_burst_packed_length_221 <= 1)) begin
            write_burst_packed_fsm_10 <= write_burst_packed_fsm_10_init;
          end 
          if(write_burst_block_ram_wvalid_217 && 0) begin
            write_burst_packed_fsm_10 <= write_burst_packed_fsm_10_init;
          end 
          if(write_burst_block_ram_wquit_218) begin
            write_burst_packed_fsm_10 <= write_burst_packed_fsm_10_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_block_fsm_11_1 = 1;
  localparam write_burst_block_fsm_11_2 = 2;
  localparam write_burst_block_fsm_11_3 = 3;
  localparam write_burst_block_fsm_11_4 = 4;
  localparam write_burst_block_fsm_11_5 = 5;
  localparam write_burst_block_fsm_11_6 = 6;
  localparam write_burst_block_fsm_11_7 = 7;
  localparam write_burst_block_fsm_11_8 = 8;
  localparam write_burst_block_fsm_11_9 = 9;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
      write_burst_block_length_231 <= 0;
      write_burst_block_blocksize_232 <= 0;
      write_burst_block_done_233 <= 0;
      write_burst_block_count_234 <= 0;
    end else begin
      case(write_burst_block_fsm_11)
        write_burst_block_fsm_11_init: begin
          write_burst_block_length_231 <= _maxi_read_local_size_buf;
          write_burst_block_blocksize_232 <= _maxi_read_local_blocksize_buf;
          write_burst_block_done_233 <= 0;
          write_burst_block_count_234 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_1;
          end 
        end
        write_burst_block_fsm_11_1: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_231 <= write_burst_block_length_231 - 1;
            write_burst_block_done_233 <= 0;
            write_burst_block_count_234 <= write_burst_block_count_234 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_231 <= 1)) begin
            write_burst_block_done_233 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_233 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_234 == write_burst_block_blocksize_232 - 1)) begin
            write_burst_block_count_234 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_234 == write_burst_block_blocksize_232 - 1)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_2;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_231 <= 1)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
          if(0) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
        end
        write_burst_block_fsm_11_2: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_231 <= write_burst_block_length_231 - 1;
            write_burst_block_done_233 <= 0;
            write_burst_block_count_234 <= write_burst_block_count_234 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_231 <= 1)) begin
            write_burst_block_done_233 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_233 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_234 == write_burst_block_blocksize_232 - 1)) begin
            write_burst_block_count_234 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_234 == write_burst_block_blocksize_232 - 1)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_3;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_231 <= 1)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
          if(0) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
        end
        write_burst_block_fsm_11_3: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_231 <= write_burst_block_length_231 - 1;
            write_burst_block_done_233 <= 0;
            write_burst_block_count_234 <= write_burst_block_count_234 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_231 <= 1)) begin
            write_burst_block_done_233 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_233 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_234 == write_burst_block_blocksize_232 - 1)) begin
            write_burst_block_count_234 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_234 == write_burst_block_blocksize_232 - 1)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_4;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_231 <= 1)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
          if(0) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
        end
        write_burst_block_fsm_11_4: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_231 <= write_burst_block_length_231 - 1;
            write_burst_block_done_233 <= 0;
            write_burst_block_count_234 <= write_burst_block_count_234 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_231 <= 1)) begin
            write_burst_block_done_233 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_233 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_234 == write_burst_block_blocksize_232 - 1)) begin
            write_burst_block_count_234 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_234 == write_burst_block_blocksize_232 - 1)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_5;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_231 <= 1)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
          if(0) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
        end
        write_burst_block_fsm_11_5: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_231 <= write_burst_block_length_231 - 1;
            write_burst_block_done_233 <= 0;
            write_burst_block_count_234 <= write_burst_block_count_234 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_231 <= 1)) begin
            write_burst_block_done_233 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_233 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_234 == write_burst_block_blocksize_232 - 1)) begin
            write_burst_block_count_234 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_234 == write_burst_block_blocksize_232 - 1)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_6;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_231 <= 1)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
          if(0) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
        end
        write_burst_block_fsm_11_6: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_231 <= write_burst_block_length_231 - 1;
            write_burst_block_done_233 <= 0;
            write_burst_block_count_234 <= write_burst_block_count_234 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_231 <= 1)) begin
            write_burst_block_done_233 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_233 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_234 == write_burst_block_blocksize_232 - 1)) begin
            write_burst_block_count_234 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_234 == write_burst_block_blocksize_232 - 1)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_7;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_231 <= 1)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
          if(0) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
        end
        write_burst_block_fsm_11_7: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_231 <= write_burst_block_length_231 - 1;
            write_burst_block_done_233 <= 0;
            write_burst_block_count_234 <= write_burst_block_count_234 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_231 <= 1)) begin
            write_burst_block_done_233 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_233 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_234 == write_burst_block_blocksize_232 - 1)) begin
            write_burst_block_count_234 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_234 == write_burst_block_blocksize_232 - 1)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_8;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_231 <= 1)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
          if(0) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
        end
        write_burst_block_fsm_11_8: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_231 <= write_burst_block_length_231 - 1;
            write_burst_block_done_233 <= 0;
            write_burst_block_count_234 <= write_burst_block_count_234 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_231 <= 1)) begin
            write_burst_block_done_233 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_233 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_234 == write_burst_block_blocksize_232 - 1)) begin
            write_burst_block_count_234 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_234 == write_burst_block_blocksize_232 - 1)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_9;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_231 <= 1)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
          if(0) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
        end
        write_burst_block_fsm_11_9: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_231 <= write_burst_block_length_231 - 1;
            write_burst_block_done_233 <= 0;
            write_burst_block_count_234 <= write_burst_block_count_234 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_231 <= 1)) begin
            write_burst_block_done_233 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_233 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_234 == write_burst_block_blocksize_232 - 1)) begin
            write_burst_block_count_234 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_234 == write_burst_block_blocksize_232 - 1)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_231 <= 1)) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
          if(0) begin
            write_burst_block_fsm_11 <= write_burst_block_fsm_11_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_12_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_12 <= write_burst_packed_fsm_12_init;
      write_burst_packed_addr_245 <= 0;
      write_burst_packed_stride_246 <= 0;
      write_burst_packed_length_247 <= 0;
      write_burst_packed_done_248 <= 0;
    end else begin
      case(write_burst_packed_fsm_12)
        write_burst_packed_fsm_12_init: begin
          write_burst_packed_addr_245 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_246 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_247 <= _maxi_read_local_size_buf;
          write_burst_packed_done_248 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 4) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_12 <= write_burst_packed_fsm_12_1;
          end 
        end
        write_burst_packed_fsm_12_1: begin
          if(write_burst_block_ram_wvalid_243) begin
            write_burst_packed_addr_245 <= write_burst_packed_addr_245 + write_burst_packed_stride_246;
            write_burst_packed_length_247 <= write_burst_packed_length_247 - 1;
            write_burst_packed_done_248 <= 0;
          end 
          if(write_burst_block_ram_wvalid_243 && (write_burst_packed_length_247 <= 1)) begin
            write_burst_packed_done_248 <= 1;
          end 
          if(write_burst_block_ram_wvalid_243 && 0) begin
            write_burst_packed_done_248 <= 1;
          end 
          if(write_burst_block_ram_wvalid_243 && (write_burst_packed_length_247 <= 1)) begin
            write_burst_packed_fsm_12 <= write_burst_packed_fsm_12_init;
          end 
          if(write_burst_block_ram_wvalid_243 && 0) begin
            write_burst_packed_fsm_12 <= write_burst_packed_fsm_12_init;
          end 
          if(write_burst_block_ram_wquit_244) begin
            write_burst_packed_fsm_12 <= write_burst_packed_fsm_12_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_13_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_13 <= write_burst_packed_fsm_13_init;
      write_burst_packed_addr_259 <= 0;
      write_burst_packed_stride_260 <= 0;
      write_burst_packed_length_261 <= 0;
      write_burst_packed_done_262 <= 0;
    end else begin
      case(write_burst_packed_fsm_13)
        write_burst_packed_fsm_13_init: begin
          write_burst_packed_addr_259 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_260 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_261 <= _maxi_read_local_size_buf;
          write_burst_packed_done_262 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 4) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_13 <= write_burst_packed_fsm_13_1;
          end 
        end
        write_burst_packed_fsm_13_1: begin
          if(write_burst_block_ram_wvalid_257) begin
            write_burst_packed_addr_259 <= write_burst_packed_addr_259 + write_burst_packed_stride_260;
            write_burst_packed_length_261 <= write_burst_packed_length_261 - 1;
            write_burst_packed_done_262 <= 0;
          end 
          if(write_burst_block_ram_wvalid_257 && (write_burst_packed_length_261 <= 1)) begin
            write_burst_packed_done_262 <= 1;
          end 
          if(write_burst_block_ram_wvalid_257 && 0) begin
            write_burst_packed_done_262 <= 1;
          end 
          if(write_burst_block_ram_wvalid_257 && (write_burst_packed_length_261 <= 1)) begin
            write_burst_packed_fsm_13 <= write_burst_packed_fsm_13_init;
          end 
          if(write_burst_block_ram_wvalid_257 && 0) begin
            write_burst_packed_fsm_13 <= write_burst_packed_fsm_13_init;
          end 
          if(write_burst_block_ram_wquit_258) begin
            write_burst_packed_fsm_13 <= write_burst_packed_fsm_13_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_14_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_14 <= write_burst_packed_fsm_14_init;
      write_burst_packed_addr_273 <= 0;
      write_burst_packed_stride_274 <= 0;
      write_burst_packed_length_275 <= 0;
      write_burst_packed_done_276 <= 0;
    end else begin
      case(write_burst_packed_fsm_14)
        write_burst_packed_fsm_14_init: begin
          write_burst_packed_addr_273 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_274 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_275 <= _maxi_read_local_size_buf;
          write_burst_packed_done_276 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 4) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_14 <= write_burst_packed_fsm_14_1;
          end 
        end
        write_burst_packed_fsm_14_1: begin
          if(write_burst_block_ram_wvalid_271) begin
            write_burst_packed_addr_273 <= write_burst_packed_addr_273 + write_burst_packed_stride_274;
            write_burst_packed_length_275 <= write_burst_packed_length_275 - 1;
            write_burst_packed_done_276 <= 0;
          end 
          if(write_burst_block_ram_wvalid_271 && (write_burst_packed_length_275 <= 1)) begin
            write_burst_packed_done_276 <= 1;
          end 
          if(write_burst_block_ram_wvalid_271 && 0) begin
            write_burst_packed_done_276 <= 1;
          end 
          if(write_burst_block_ram_wvalid_271 && (write_burst_packed_length_275 <= 1)) begin
            write_burst_packed_fsm_14 <= write_burst_packed_fsm_14_init;
          end 
          if(write_burst_block_ram_wvalid_271 && 0) begin
            write_burst_packed_fsm_14 <= write_burst_packed_fsm_14_init;
          end 
          if(write_burst_block_ram_wquit_272) begin
            write_burst_packed_fsm_14 <= write_burst_packed_fsm_14_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_block_fsm_15_1 = 1;
  localparam write_burst_block_fsm_15_2 = 2;
  localparam write_burst_block_fsm_15_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_block_fsm_15 <= write_burst_block_fsm_15_init;
      write_burst_block_length_285 <= 0;
      write_burst_block_blocksize_286 <= 0;
      write_burst_block_done_287 <= 0;
      write_burst_block_count_288 <= 0;
    end else begin
      case(write_burst_block_fsm_15)
        write_burst_block_fsm_15_init: begin
          write_burst_block_length_285 <= _maxi_read_local_size_buf;
          write_burst_block_blocksize_286 <= _maxi_read_local_blocksize_buf;
          write_burst_block_done_287 <= 0;
          write_burst_block_count_288 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 4) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_block_fsm_15 <= write_burst_block_fsm_15_1;
          end 
        end
        write_burst_block_fsm_15_1: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_285 <= write_burst_block_length_285 - 1;
            write_burst_block_done_287 <= 0;
            write_burst_block_count_288 <= write_burst_block_count_288 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_285 <= 1)) begin
            write_burst_block_done_287 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_287 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_288 == write_burst_block_blocksize_286 - 1)) begin
            write_burst_block_count_288 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_288 == write_burst_block_blocksize_286 - 1)) begin
            write_burst_block_fsm_15 <= write_burst_block_fsm_15_2;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_285 <= 1)) begin
            write_burst_block_fsm_15 <= write_burst_block_fsm_15_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_15 <= write_burst_block_fsm_15_init;
          end 
          if(0) begin
            write_burst_block_fsm_15 <= write_burst_block_fsm_15_init;
          end 
        end
        write_burst_block_fsm_15_2: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_285 <= write_burst_block_length_285 - 1;
            write_burst_block_done_287 <= 0;
            write_burst_block_count_288 <= write_burst_block_count_288 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_285 <= 1)) begin
            write_burst_block_done_287 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_287 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_288 == write_burst_block_blocksize_286 - 1)) begin
            write_burst_block_count_288 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_288 == write_burst_block_blocksize_286 - 1)) begin
            write_burst_block_fsm_15 <= write_burst_block_fsm_15_3;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_285 <= 1)) begin
            write_burst_block_fsm_15 <= write_burst_block_fsm_15_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_15 <= write_burst_block_fsm_15_init;
          end 
          if(0) begin
            write_burst_block_fsm_15 <= write_burst_block_fsm_15_init;
          end 
        end
        write_burst_block_fsm_15_3: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_285 <= write_burst_block_length_285 - 1;
            write_burst_block_done_287 <= 0;
            write_burst_block_count_288 <= write_burst_block_count_288 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_285 <= 1)) begin
            write_burst_block_done_287 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_287 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_288 == write_burst_block_blocksize_286 - 1)) begin
            write_burst_block_count_288 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_288 == write_burst_block_blocksize_286 - 1)) begin
            write_burst_block_fsm_15 <= write_burst_block_fsm_15_1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_285 <= 1)) begin
            write_burst_block_fsm_15 <= write_burst_block_fsm_15_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_15 <= write_burst_block_fsm_15_init;
          end 
          if(0) begin
            write_burst_block_fsm_15 <= write_burst_block_fsm_15_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_16_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_16 <= write_burst_packed_fsm_16_init;
      write_burst_packed_addr_299 <= 0;
      write_burst_packed_stride_300 <= 0;
      write_burst_packed_length_301 <= 0;
      write_burst_packed_done_302 <= 0;
    end else begin
      case(write_burst_packed_fsm_16)
        write_burst_packed_fsm_16_init: begin
          write_burst_packed_addr_299 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_300 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_301 <= _maxi_read_local_size_buf;
          write_burst_packed_done_302 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 5) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_16 <= write_burst_packed_fsm_16_1;
          end 
        end
        write_burst_packed_fsm_16_1: begin
          if(write_burst_block_ram_wvalid_297) begin
            write_burst_packed_addr_299 <= write_burst_packed_addr_299 + write_burst_packed_stride_300;
            write_burst_packed_length_301 <= write_burst_packed_length_301 - 1;
            write_burst_packed_done_302 <= 0;
          end 
          if(write_burst_block_ram_wvalid_297 && (write_burst_packed_length_301 <= 1)) begin
            write_burst_packed_done_302 <= 1;
          end 
          if(write_burst_block_ram_wvalid_297 && 0) begin
            write_burst_packed_done_302 <= 1;
          end 
          if(write_burst_block_ram_wvalid_297 && (write_burst_packed_length_301 <= 1)) begin
            write_burst_packed_fsm_16 <= write_burst_packed_fsm_16_init;
          end 
          if(write_burst_block_ram_wvalid_297 && 0) begin
            write_burst_packed_fsm_16 <= write_burst_packed_fsm_16_init;
          end 
          if(write_burst_block_ram_wquit_298) begin
            write_burst_packed_fsm_16 <= write_burst_packed_fsm_16_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_17_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_17 <= write_burst_packed_fsm_17_init;
      write_burst_packed_addr_313 <= 0;
      write_burst_packed_stride_314 <= 0;
      write_burst_packed_length_315 <= 0;
      write_burst_packed_done_316 <= 0;
    end else begin
      case(write_burst_packed_fsm_17)
        write_burst_packed_fsm_17_init: begin
          write_burst_packed_addr_313 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_314 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_315 <= _maxi_read_local_size_buf;
          write_burst_packed_done_316 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 5) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_17 <= write_burst_packed_fsm_17_1;
          end 
        end
        write_burst_packed_fsm_17_1: begin
          if(write_burst_block_ram_wvalid_311) begin
            write_burst_packed_addr_313 <= write_burst_packed_addr_313 + write_burst_packed_stride_314;
            write_burst_packed_length_315 <= write_burst_packed_length_315 - 1;
            write_burst_packed_done_316 <= 0;
          end 
          if(write_burst_block_ram_wvalid_311 && (write_burst_packed_length_315 <= 1)) begin
            write_burst_packed_done_316 <= 1;
          end 
          if(write_burst_block_ram_wvalid_311 && 0) begin
            write_burst_packed_done_316 <= 1;
          end 
          if(write_burst_block_ram_wvalid_311 && (write_burst_packed_length_315 <= 1)) begin
            write_burst_packed_fsm_17 <= write_burst_packed_fsm_17_init;
          end 
          if(write_burst_block_ram_wvalid_311 && 0) begin
            write_burst_packed_fsm_17 <= write_burst_packed_fsm_17_init;
          end 
          if(write_burst_block_ram_wquit_312) begin
            write_burst_packed_fsm_17 <= write_burst_packed_fsm_17_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_18_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_18 <= write_burst_packed_fsm_18_init;
      write_burst_packed_addr_327 <= 0;
      write_burst_packed_stride_328 <= 0;
      write_burst_packed_length_329 <= 0;
      write_burst_packed_done_330 <= 0;
    end else begin
      case(write_burst_packed_fsm_18)
        write_burst_packed_fsm_18_init: begin
          write_burst_packed_addr_327 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_328 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_329 <= _maxi_read_local_size_buf;
          write_burst_packed_done_330 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 5) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_18 <= write_burst_packed_fsm_18_1;
          end 
        end
        write_burst_packed_fsm_18_1: begin
          if(write_burst_block_ram_wvalid_325) begin
            write_burst_packed_addr_327 <= write_burst_packed_addr_327 + write_burst_packed_stride_328;
            write_burst_packed_length_329 <= write_burst_packed_length_329 - 1;
            write_burst_packed_done_330 <= 0;
          end 
          if(write_burst_block_ram_wvalid_325 && (write_burst_packed_length_329 <= 1)) begin
            write_burst_packed_done_330 <= 1;
          end 
          if(write_burst_block_ram_wvalid_325 && 0) begin
            write_burst_packed_done_330 <= 1;
          end 
          if(write_burst_block_ram_wvalid_325 && (write_burst_packed_length_329 <= 1)) begin
            write_burst_packed_fsm_18 <= write_burst_packed_fsm_18_init;
          end 
          if(write_burst_block_ram_wvalid_325 && 0) begin
            write_burst_packed_fsm_18 <= write_burst_packed_fsm_18_init;
          end 
          if(write_burst_block_ram_wquit_326) begin
            write_burst_packed_fsm_18 <= write_burst_packed_fsm_18_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_block_fsm_19_1 = 1;
  localparam write_burst_block_fsm_19_2 = 2;
  localparam write_burst_block_fsm_19_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_block_fsm_19 <= write_burst_block_fsm_19_init;
      write_burst_block_length_339 <= 0;
      write_burst_block_blocksize_340 <= 0;
      write_burst_block_done_341 <= 0;
      write_burst_block_count_342 <= 0;
    end else begin
      case(write_burst_block_fsm_19)
        write_burst_block_fsm_19_init: begin
          write_burst_block_length_339 <= _maxi_read_local_size_buf;
          write_burst_block_blocksize_340 <= _maxi_read_local_blocksize_buf;
          write_burst_block_done_341 <= 0;
          write_burst_block_count_342 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 5) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_block_fsm_19 <= write_burst_block_fsm_19_1;
          end 
        end
        write_burst_block_fsm_19_1: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_339 <= write_burst_block_length_339 - 1;
            write_burst_block_done_341 <= 0;
            write_burst_block_count_342 <= write_burst_block_count_342 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_339 <= 1)) begin
            write_burst_block_done_341 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_341 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_342 == write_burst_block_blocksize_340 - 1)) begin
            write_burst_block_count_342 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_342 == write_burst_block_blocksize_340 - 1)) begin
            write_burst_block_fsm_19 <= write_burst_block_fsm_19_2;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_339 <= 1)) begin
            write_burst_block_fsm_19 <= write_burst_block_fsm_19_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_19 <= write_burst_block_fsm_19_init;
          end 
          if(0) begin
            write_burst_block_fsm_19 <= write_burst_block_fsm_19_init;
          end 
        end
        write_burst_block_fsm_19_2: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_339 <= write_burst_block_length_339 - 1;
            write_burst_block_done_341 <= 0;
            write_burst_block_count_342 <= write_burst_block_count_342 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_339 <= 1)) begin
            write_burst_block_done_341 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_341 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_342 == write_burst_block_blocksize_340 - 1)) begin
            write_burst_block_count_342 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_342 == write_burst_block_blocksize_340 - 1)) begin
            write_burst_block_fsm_19 <= write_burst_block_fsm_19_3;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_339 <= 1)) begin
            write_burst_block_fsm_19 <= write_burst_block_fsm_19_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_19 <= write_burst_block_fsm_19_init;
          end 
          if(0) begin
            write_burst_block_fsm_19 <= write_burst_block_fsm_19_init;
          end 
        end
        write_burst_block_fsm_19_3: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_339 <= write_burst_block_length_339 - 1;
            write_burst_block_done_341 <= 0;
            write_burst_block_count_342 <= write_burst_block_count_342 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_339 <= 1)) begin
            write_burst_block_done_341 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_341 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_342 == write_burst_block_blocksize_340 - 1)) begin
            write_burst_block_count_342 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_342 == write_burst_block_blocksize_340 - 1)) begin
            write_burst_block_fsm_19 <= write_burst_block_fsm_19_1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_339 <= 1)) begin
            write_burst_block_fsm_19 <= write_burst_block_fsm_19_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_19 <= write_burst_block_fsm_19_init;
          end 
          if(0) begin
            write_burst_block_fsm_19 <= write_burst_block_fsm_19_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_20_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_20 <= write_burst_packed_fsm_20_init;
      write_burst_packed_addr_353 <= 0;
      write_burst_packed_stride_354 <= 0;
      write_burst_packed_length_355 <= 0;
      write_burst_packed_done_356 <= 0;
    end else begin
      case(write_burst_packed_fsm_20)
        write_burst_packed_fsm_20_init: begin
          write_burst_packed_addr_353 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_354 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_355 <= _maxi_read_local_size_buf;
          write_burst_packed_done_356 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 6) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_20 <= write_burst_packed_fsm_20_1;
          end 
        end
        write_burst_packed_fsm_20_1: begin
          if(write_burst_block_ram_wvalid_351) begin
            write_burst_packed_addr_353 <= write_burst_packed_addr_353 + write_burst_packed_stride_354;
            write_burst_packed_length_355 <= write_burst_packed_length_355 - 1;
            write_burst_packed_done_356 <= 0;
          end 
          if(write_burst_block_ram_wvalid_351 && (write_burst_packed_length_355 <= 1)) begin
            write_burst_packed_done_356 <= 1;
          end 
          if(write_burst_block_ram_wvalid_351 && 0) begin
            write_burst_packed_done_356 <= 1;
          end 
          if(write_burst_block_ram_wvalid_351 && (write_burst_packed_length_355 <= 1)) begin
            write_burst_packed_fsm_20 <= write_burst_packed_fsm_20_init;
          end 
          if(write_burst_block_ram_wvalid_351 && 0) begin
            write_burst_packed_fsm_20 <= write_burst_packed_fsm_20_init;
          end 
          if(write_burst_block_ram_wquit_352) begin
            write_burst_packed_fsm_20 <= write_burst_packed_fsm_20_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_21_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_21 <= write_burst_packed_fsm_21_init;
      write_burst_packed_addr_367 <= 0;
      write_burst_packed_stride_368 <= 0;
      write_burst_packed_length_369 <= 0;
      write_burst_packed_done_370 <= 0;
    end else begin
      case(write_burst_packed_fsm_21)
        write_burst_packed_fsm_21_init: begin
          write_burst_packed_addr_367 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_368 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_369 <= _maxi_read_local_size_buf;
          write_burst_packed_done_370 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 6) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_21 <= write_burst_packed_fsm_21_1;
          end 
        end
        write_burst_packed_fsm_21_1: begin
          if(write_burst_block_ram_wvalid_365) begin
            write_burst_packed_addr_367 <= write_burst_packed_addr_367 + write_burst_packed_stride_368;
            write_burst_packed_length_369 <= write_burst_packed_length_369 - 1;
            write_burst_packed_done_370 <= 0;
          end 
          if(write_burst_block_ram_wvalid_365 && (write_burst_packed_length_369 <= 1)) begin
            write_burst_packed_done_370 <= 1;
          end 
          if(write_burst_block_ram_wvalid_365 && 0) begin
            write_burst_packed_done_370 <= 1;
          end 
          if(write_burst_block_ram_wvalid_365 && (write_burst_packed_length_369 <= 1)) begin
            write_burst_packed_fsm_21 <= write_burst_packed_fsm_21_init;
          end 
          if(write_burst_block_ram_wvalid_365 && 0) begin
            write_burst_packed_fsm_21 <= write_burst_packed_fsm_21_init;
          end 
          if(write_burst_block_ram_wquit_366) begin
            write_burst_packed_fsm_21 <= write_burst_packed_fsm_21_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_22_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_22 <= write_burst_packed_fsm_22_init;
      write_burst_packed_addr_381 <= 0;
      write_burst_packed_stride_382 <= 0;
      write_burst_packed_length_383 <= 0;
      write_burst_packed_done_384 <= 0;
    end else begin
      case(write_burst_packed_fsm_22)
        write_burst_packed_fsm_22_init: begin
          write_burst_packed_addr_381 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_382 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_383 <= _maxi_read_local_size_buf;
          write_burst_packed_done_384 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 6) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_22 <= write_burst_packed_fsm_22_1;
          end 
        end
        write_burst_packed_fsm_22_1: begin
          if(write_burst_block_ram_wvalid_379) begin
            write_burst_packed_addr_381 <= write_burst_packed_addr_381 + write_burst_packed_stride_382;
            write_burst_packed_length_383 <= write_burst_packed_length_383 - 1;
            write_burst_packed_done_384 <= 0;
          end 
          if(write_burst_block_ram_wvalid_379 && (write_burst_packed_length_383 <= 1)) begin
            write_burst_packed_done_384 <= 1;
          end 
          if(write_burst_block_ram_wvalid_379 && 0) begin
            write_burst_packed_done_384 <= 1;
          end 
          if(write_burst_block_ram_wvalid_379 && (write_burst_packed_length_383 <= 1)) begin
            write_burst_packed_fsm_22 <= write_burst_packed_fsm_22_init;
          end 
          if(write_burst_block_ram_wvalid_379 && 0) begin
            write_burst_packed_fsm_22 <= write_burst_packed_fsm_22_init;
          end 
          if(write_burst_block_ram_wquit_380) begin
            write_burst_packed_fsm_22 <= write_burst_packed_fsm_22_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_block_fsm_23_1 = 1;
  localparam write_burst_block_fsm_23_2 = 2;
  localparam write_burst_block_fsm_23_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_block_fsm_23 <= write_burst_block_fsm_23_init;
      write_burst_block_length_393 <= 0;
      write_burst_block_blocksize_394 <= 0;
      write_burst_block_done_395 <= 0;
      write_burst_block_count_396 <= 0;
    end else begin
      case(write_burst_block_fsm_23)
        write_burst_block_fsm_23_init: begin
          write_burst_block_length_393 <= _maxi_read_local_size_buf;
          write_burst_block_blocksize_394 <= _maxi_read_local_blocksize_buf;
          write_burst_block_done_395 <= 0;
          write_burst_block_count_396 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 6) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_block_fsm_23 <= write_burst_block_fsm_23_1;
          end 
        end
        write_burst_block_fsm_23_1: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_393 <= write_burst_block_length_393 - 1;
            write_burst_block_done_395 <= 0;
            write_burst_block_count_396 <= write_burst_block_count_396 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_393 <= 1)) begin
            write_burst_block_done_395 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_395 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_396 == write_burst_block_blocksize_394 - 1)) begin
            write_burst_block_count_396 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_396 == write_burst_block_blocksize_394 - 1)) begin
            write_burst_block_fsm_23 <= write_burst_block_fsm_23_2;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_393 <= 1)) begin
            write_burst_block_fsm_23 <= write_burst_block_fsm_23_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_23 <= write_burst_block_fsm_23_init;
          end 
          if(0) begin
            write_burst_block_fsm_23 <= write_burst_block_fsm_23_init;
          end 
        end
        write_burst_block_fsm_23_2: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_393 <= write_burst_block_length_393 - 1;
            write_burst_block_done_395 <= 0;
            write_burst_block_count_396 <= write_burst_block_count_396 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_393 <= 1)) begin
            write_burst_block_done_395 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_395 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_396 == write_burst_block_blocksize_394 - 1)) begin
            write_burst_block_count_396 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_396 == write_burst_block_blocksize_394 - 1)) begin
            write_burst_block_fsm_23 <= write_burst_block_fsm_23_3;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_393 <= 1)) begin
            write_burst_block_fsm_23 <= write_burst_block_fsm_23_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_23 <= write_burst_block_fsm_23_init;
          end 
          if(0) begin
            write_burst_block_fsm_23 <= write_burst_block_fsm_23_init;
          end 
        end
        write_burst_block_fsm_23_3: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_393 <= write_burst_block_length_393 - 1;
            write_burst_block_done_395 <= 0;
            write_burst_block_count_396 <= write_burst_block_count_396 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_393 <= 1)) begin
            write_burst_block_done_395 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_395 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_396 == write_burst_block_blocksize_394 - 1)) begin
            write_burst_block_count_396 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_396 == write_burst_block_blocksize_394 - 1)) begin
            write_burst_block_fsm_23 <= write_burst_block_fsm_23_1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_393 <= 1)) begin
            write_burst_block_fsm_23 <= write_burst_block_fsm_23_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_23 <= write_burst_block_fsm_23_init;
          end 
          if(0) begin
            write_burst_block_fsm_23 <= write_burst_block_fsm_23_init;
          end 
        end
      endcase
    end
  end

  localparam conv2d_24_comp_fsm_1 = 1;
  localparam conv2d_24_comp_fsm_2 = 2;
  localparam conv2d_24_comp_fsm_3 = 3;
  localparam conv2d_24_comp_fsm_4 = 4;
  localparam conv2d_24_comp_fsm_5 = 5;
  localparam conv2d_24_comp_fsm_6 = 6;

  always @(posedge CLK) begin
    if(RST) begin
      conv2d_24_comp_fsm <= conv2d_24_comp_fsm_init;
      conv2d_24_stream_act_local_0 <= 0;
      conv2d_24_stream_act_local_1 <= 0;
      conv2d_24_stream_act_local_2 <= 0;
      conv2d_24_stream_act_local_3 <= 0;
      conv2d_24_stream_act_local_4 <= 0;
      conv2d_24_stream_act_local_5 <= 0;
      conv2d_24_stream_act_local_6 <= 0;
      conv2d_24_stream_act_local_7 <= 0;
      conv2d_24_stream_act_local_8 <= 0;
      conv2d_24_stream_out_local_col <= 0;
      conv2d_24_stream_out_local_val <= 0;
      conv2d_24_col_count <= 0;
      conv2d_24_col_select <= 0;
      conv2d_24_filter_page_comp_offset_buf <= 0;
      conv2d_24_act_page_comp_offset_buf_0 <= 0;
      conv2d_24_act_page_comp_offset_buf_1 <= 0;
      conv2d_24_act_page_comp_offset_buf_2 <= 0;
      conv2d_24_out_page_comp_offset_buf <= 0;
      conv2d_24_row_count_buf <= 0;
      conv2d_24_row_select_buf <= 0;
      conv2d_24_och_count_buf <= 0;
      conv2d_24_next_stream_num_ops <= 0;
      conv2d_24_stream_pad_masks <= 0;
      conv2d_24_sync_comp_count <= 0;
    end else begin
      if(_stream_conv2d_24_sink_stop) begin
        conv2d_24_sync_comp_count <= conv2d_24_sync_comp_count + 1;
      end 
      if(control_conv2d_24 == 6) begin
        conv2d_24_sync_comp_count <= 0;
      end 
      case(conv2d_24_comp_fsm)
        conv2d_24_comp_fsm_init: begin
          if((control_conv2d_24 == 25) && !conv2d_24_skip_comp) begin
            conv2d_24_comp_fsm <= conv2d_24_comp_fsm_1;
          end 
        end
        conv2d_24_comp_fsm_1: begin
          conv2d_24_stream_act_local_0 <= 0;
          if(cparam_conv2d_24_stream_act_local_small_flags_0) begin
            conv2d_24_stream_act_local_0 <= cparam_conv2d_24_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_24_stream_act_local_large_flags_0) begin
            conv2d_24_stream_act_local_0 <= cparam_conv2d_24_stream_act_local_large_offset;
          end 
          conv2d_24_stream_act_local_1 <= 0;
          if(cparam_conv2d_24_stream_act_local_small_flags_1) begin
            conv2d_24_stream_act_local_1 <= cparam_conv2d_24_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_24_stream_act_local_large_flags_1) begin
            conv2d_24_stream_act_local_1 <= cparam_conv2d_24_stream_act_local_large_offset;
          end 
          conv2d_24_stream_act_local_2 <= 0;
          if(cparam_conv2d_24_stream_act_local_small_flags_2) begin
            conv2d_24_stream_act_local_2 <= cparam_conv2d_24_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_24_stream_act_local_large_flags_2) begin
            conv2d_24_stream_act_local_2 <= cparam_conv2d_24_stream_act_local_large_offset;
          end 
          conv2d_24_stream_act_local_3 <= 0;
          if(cparam_conv2d_24_stream_act_local_small_flags_0) begin
            conv2d_24_stream_act_local_3 <= cparam_conv2d_24_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_24_stream_act_local_large_flags_0) begin
            conv2d_24_stream_act_local_3 <= cparam_conv2d_24_stream_act_local_large_offset;
          end 
          conv2d_24_stream_act_local_4 <= 0;
          if(cparam_conv2d_24_stream_act_local_small_flags_1) begin
            conv2d_24_stream_act_local_4 <= cparam_conv2d_24_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_24_stream_act_local_large_flags_1) begin
            conv2d_24_stream_act_local_4 <= cparam_conv2d_24_stream_act_local_large_offset;
          end 
          conv2d_24_stream_act_local_5 <= 0;
          if(cparam_conv2d_24_stream_act_local_small_flags_2) begin
            conv2d_24_stream_act_local_5 <= cparam_conv2d_24_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_24_stream_act_local_large_flags_2) begin
            conv2d_24_stream_act_local_5 <= cparam_conv2d_24_stream_act_local_large_offset;
          end 
          conv2d_24_stream_act_local_6 <= 0;
          if(cparam_conv2d_24_stream_act_local_small_flags_0) begin
            conv2d_24_stream_act_local_6 <= cparam_conv2d_24_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_24_stream_act_local_large_flags_0) begin
            conv2d_24_stream_act_local_6 <= cparam_conv2d_24_stream_act_local_large_offset;
          end 
          conv2d_24_stream_act_local_7 <= 0;
          if(cparam_conv2d_24_stream_act_local_small_flags_1) begin
            conv2d_24_stream_act_local_7 <= cparam_conv2d_24_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_24_stream_act_local_large_flags_1) begin
            conv2d_24_stream_act_local_7 <= cparam_conv2d_24_stream_act_local_large_offset;
          end 
          conv2d_24_stream_act_local_8 <= 0;
          if(cparam_conv2d_24_stream_act_local_small_flags_2) begin
            conv2d_24_stream_act_local_8 <= cparam_conv2d_24_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_24_stream_act_local_large_flags_2) begin
            conv2d_24_stream_act_local_8 <= cparam_conv2d_24_stream_act_local_large_offset;
          end 
          conv2d_24_stream_out_local_col <= 0;
          if((cparam_conv2d_24_data_stationary == 1) && (conv2d_24_och_count == 0)) begin
            conv2d_24_stream_out_local_val <= 0;
          end 
          conv2d_24_col_count <= 0;
          conv2d_24_col_select <= cparam_conv2d_24_col_select_initval;
          conv2d_24_filter_page_comp_offset_buf <= conv2d_24_filter_page_comp_offset;
          conv2d_24_act_page_comp_offset_buf_0 <= conv2d_24_act_page_comp_offset_0;
          conv2d_24_act_page_comp_offset_buf_1 <= conv2d_24_act_page_comp_offset_1;
          conv2d_24_act_page_comp_offset_buf_2 <= conv2d_24_act_page_comp_offset_2;
          conv2d_24_out_page_comp_offset_buf <= conv2d_24_out_page_comp_offset;
          conv2d_24_row_count_buf <= conv2d_24_row_count;
          conv2d_24_row_select_buf <= conv2d_24_row_select;
          conv2d_24_och_count_buf <= conv2d_24_och_count;
          conv2d_24_next_stream_num_ops <= (conv2d_24_och_count >= cparam_conv2d_24_max_och_count)? cparam_conv2d_24_stream_num_ops_res : cparam_conv2d_24_stream_num_ops;
          conv2d_24_comp_fsm <= conv2d_24_comp_fsm_2;
        end
        conv2d_24_comp_fsm_2: begin
          conv2d_24_stream_pad_masks <= { conv2d_24_stream_pad_mask_2_2, conv2d_24_stream_pad_mask_2_1, conv2d_24_stream_pad_mask_2_0, conv2d_24_stream_pad_mask_1_2, conv2d_24_stream_pad_mask_1_1, conv2d_24_stream_pad_mask_1_0, conv2d_24_stream_pad_mask_0_2, conv2d_24_stream_pad_mask_0_1, conv2d_24_stream_pad_mask_0_0 };
          conv2d_24_comp_fsm <= conv2d_24_comp_fsm_3;
        end
        conv2d_24_comp_fsm_3: begin
          conv2d_24_comp_fsm <= conv2d_24_comp_fsm_4;
          conv2d_24_comp_fsm <= conv2d_24_comp_fsm_4;
          conv2d_24_comp_fsm <= conv2d_24_comp_fsm_4;
          conv2d_24_comp_fsm <= conv2d_24_comp_fsm_4;
          conv2d_24_comp_fsm <= conv2d_24_comp_fsm_4;
          conv2d_24_comp_fsm <= conv2d_24_comp_fsm_4;
          conv2d_24_comp_fsm <= conv2d_24_comp_fsm_4;
          conv2d_24_comp_fsm <= conv2d_24_comp_fsm_4;
          conv2d_24_comp_fsm <= conv2d_24_comp_fsm_4;
          conv2d_24_comp_fsm <= conv2d_24_comp_fsm_4;
          conv2d_24_comp_fsm <= conv2d_24_comp_fsm_4;
          conv2d_24_comp_fsm <= conv2d_24_comp_fsm_4;
          conv2d_24_comp_fsm <= conv2d_24_comp_fsm_4;
          conv2d_24_comp_fsm <= conv2d_24_comp_fsm_4;
          conv2d_24_comp_fsm <= conv2d_24_comp_fsm_4;
          conv2d_24_comp_fsm <= conv2d_24_comp_fsm_4;
          conv2d_24_comp_fsm <= conv2d_24_comp_fsm_4;
          conv2d_24_comp_fsm <= conv2d_24_comp_fsm_4;
          conv2d_24_comp_fsm <= conv2d_24_comp_fsm_4;
          conv2d_24_comp_fsm <= conv2d_24_comp_fsm_4;
          conv2d_24_comp_fsm <= conv2d_24_comp_fsm_4;
          conv2d_24_comp_fsm <= conv2d_24_comp_fsm_4;
          conv2d_24_comp_fsm <= conv2d_24_comp_fsm_4;
          conv2d_24_comp_fsm <= conv2d_24_comp_fsm_4;
          conv2d_24_comp_fsm <= conv2d_24_comp_fsm_4;
          conv2d_24_comp_fsm <= conv2d_24_comp_fsm_4;
          conv2d_24_comp_fsm <= conv2d_24_comp_fsm_4;
          conv2d_24_comp_fsm <= conv2d_24_comp_fsm_4;
          conv2d_24_comp_fsm <= conv2d_24_comp_fsm_4;
          conv2d_24_comp_fsm <= conv2d_24_comp_fsm_4;
          conv2d_24_comp_fsm <= conv2d_24_comp_fsm_4;
          conv2d_24_comp_fsm <= conv2d_24_comp_fsm_4;
          conv2d_24_comp_fsm <= conv2d_24_comp_fsm_4;
          conv2d_24_comp_fsm <= conv2d_24_comp_fsm_4;
          conv2d_24_comp_fsm <= conv2d_24_comp_fsm_4;
          conv2d_24_comp_fsm <= conv2d_24_comp_fsm_4;
          conv2d_24_comp_fsm <= conv2d_24_comp_fsm_4;
          if(_stream_conv2d_24_stream_oready) begin
            conv2d_24_comp_fsm <= conv2d_24_comp_fsm_4;
          end 
          conv2d_24_comp_fsm <= conv2d_24_comp_fsm_4;
        end
        conv2d_24_comp_fsm_4: begin
          if(!_stream_conv2d_24_source_busy) begin
            conv2d_24_comp_fsm <= conv2d_24_comp_fsm_5;
          end 
        end
        conv2d_24_comp_fsm_5: begin
          if(_stream_conv2d_24_busy) begin
            conv2d_24_comp_fsm <= conv2d_24_comp_fsm_6;
          end 
        end
        conv2d_24_comp_fsm_6: begin
          if(!((conv2d_24_col_select == 0)? cparam_conv2d_24_inc_act_laddr_conds_0 : 
          (conv2d_24_col_select == 1)? cparam_conv2d_24_inc_act_laddr_conds_1 : 
          (conv2d_24_col_select == 2)? cparam_conv2d_24_inc_act_laddr_conds_2 : 0)) begin
            conv2d_24_stream_act_local_0 <= conv2d_24_stream_act_local_0 + cparam_conv2d_24_inc_act_laddr_small;
          end 
          if((conv2d_24_col_select == 0)? cparam_conv2d_24_inc_act_laddr_conds_0 : 
          (conv2d_24_col_select == 1)? cparam_conv2d_24_inc_act_laddr_conds_1 : 
          (conv2d_24_col_select == 2)? cparam_conv2d_24_inc_act_laddr_conds_2 : 0) begin
            conv2d_24_stream_act_local_0 <= conv2d_24_stream_act_local_0 + cparam_conv2d_24_inc_act_laddr_large;
          end 
          if(conv2d_24_col_count >= cparam_conv2d_24_max_col_count) begin
            conv2d_24_stream_act_local_0 <= 0;
          end 
          if((conv2d_24_col_count >= cparam_conv2d_24_max_col_count) && cparam_conv2d_24_stream_act_local_small_flags_0) begin
            conv2d_24_stream_act_local_0 <= cparam_conv2d_24_stream_act_local_small_offset;
          end 
          if((conv2d_24_col_count >= cparam_conv2d_24_max_col_count) && cparam_conv2d_24_stream_act_local_large_flags_0) begin
            conv2d_24_stream_act_local_0 <= cparam_conv2d_24_stream_act_local_large_offset;
          end 
          if(!((conv2d_24_col_select == 0)? cparam_conv2d_24_inc_act_laddr_conds_3 : 
          (conv2d_24_col_select == 1)? cparam_conv2d_24_inc_act_laddr_conds_4 : 
          (conv2d_24_col_select == 2)? cparam_conv2d_24_inc_act_laddr_conds_5 : 0)) begin
            conv2d_24_stream_act_local_1 <= conv2d_24_stream_act_local_1 + cparam_conv2d_24_inc_act_laddr_small;
          end 
          if((conv2d_24_col_select == 0)? cparam_conv2d_24_inc_act_laddr_conds_3 : 
          (conv2d_24_col_select == 1)? cparam_conv2d_24_inc_act_laddr_conds_4 : 
          (conv2d_24_col_select == 2)? cparam_conv2d_24_inc_act_laddr_conds_5 : 0) begin
            conv2d_24_stream_act_local_1 <= conv2d_24_stream_act_local_1 + cparam_conv2d_24_inc_act_laddr_large;
          end 
          if(conv2d_24_col_count >= cparam_conv2d_24_max_col_count) begin
            conv2d_24_stream_act_local_1 <= 0;
          end 
          if((conv2d_24_col_count >= cparam_conv2d_24_max_col_count) && cparam_conv2d_24_stream_act_local_small_flags_1) begin
            conv2d_24_stream_act_local_1 <= cparam_conv2d_24_stream_act_local_small_offset;
          end 
          if((conv2d_24_col_count >= cparam_conv2d_24_max_col_count) && cparam_conv2d_24_stream_act_local_large_flags_1) begin
            conv2d_24_stream_act_local_1 <= cparam_conv2d_24_stream_act_local_large_offset;
          end 
          if(!((conv2d_24_col_select == 0)? cparam_conv2d_24_inc_act_laddr_conds_6 : 
          (conv2d_24_col_select == 1)? cparam_conv2d_24_inc_act_laddr_conds_7 : 
          (conv2d_24_col_select == 2)? cparam_conv2d_24_inc_act_laddr_conds_8 : 0)) begin
            conv2d_24_stream_act_local_2 <= conv2d_24_stream_act_local_2 + cparam_conv2d_24_inc_act_laddr_small;
          end 
          if((conv2d_24_col_select == 0)? cparam_conv2d_24_inc_act_laddr_conds_6 : 
          (conv2d_24_col_select == 1)? cparam_conv2d_24_inc_act_laddr_conds_7 : 
          (conv2d_24_col_select == 2)? cparam_conv2d_24_inc_act_laddr_conds_8 : 0) begin
            conv2d_24_stream_act_local_2 <= conv2d_24_stream_act_local_2 + cparam_conv2d_24_inc_act_laddr_large;
          end 
          if(conv2d_24_col_count >= cparam_conv2d_24_max_col_count) begin
            conv2d_24_stream_act_local_2 <= 0;
          end 
          if((conv2d_24_col_count >= cparam_conv2d_24_max_col_count) && cparam_conv2d_24_stream_act_local_small_flags_2) begin
            conv2d_24_stream_act_local_2 <= cparam_conv2d_24_stream_act_local_small_offset;
          end 
          if((conv2d_24_col_count >= cparam_conv2d_24_max_col_count) && cparam_conv2d_24_stream_act_local_large_flags_2) begin
            conv2d_24_stream_act_local_2 <= cparam_conv2d_24_stream_act_local_large_offset;
          end 
          if(!((conv2d_24_col_select == 0)? cparam_conv2d_24_inc_act_laddr_conds_9 : 
          (conv2d_24_col_select == 1)? cparam_conv2d_24_inc_act_laddr_conds_10 : 
          (conv2d_24_col_select == 2)? cparam_conv2d_24_inc_act_laddr_conds_11 : 0)) begin
            conv2d_24_stream_act_local_3 <= conv2d_24_stream_act_local_3 + cparam_conv2d_24_inc_act_laddr_small;
          end 
          if((conv2d_24_col_select == 0)? cparam_conv2d_24_inc_act_laddr_conds_9 : 
          (conv2d_24_col_select == 1)? cparam_conv2d_24_inc_act_laddr_conds_10 : 
          (conv2d_24_col_select == 2)? cparam_conv2d_24_inc_act_laddr_conds_11 : 0) begin
            conv2d_24_stream_act_local_3 <= conv2d_24_stream_act_local_3 + cparam_conv2d_24_inc_act_laddr_large;
          end 
          if(conv2d_24_col_count >= cparam_conv2d_24_max_col_count) begin
            conv2d_24_stream_act_local_3 <= 0;
          end 
          if((conv2d_24_col_count >= cparam_conv2d_24_max_col_count) && cparam_conv2d_24_stream_act_local_small_flags_0) begin
            conv2d_24_stream_act_local_3 <= cparam_conv2d_24_stream_act_local_small_offset;
          end 
          if((conv2d_24_col_count >= cparam_conv2d_24_max_col_count) && cparam_conv2d_24_stream_act_local_large_flags_0) begin
            conv2d_24_stream_act_local_3 <= cparam_conv2d_24_stream_act_local_large_offset;
          end 
          if(!((conv2d_24_col_select == 0)? cparam_conv2d_24_inc_act_laddr_conds_12 : 
          (conv2d_24_col_select == 1)? cparam_conv2d_24_inc_act_laddr_conds_13 : 
          (conv2d_24_col_select == 2)? cparam_conv2d_24_inc_act_laddr_conds_14 : 0)) begin
            conv2d_24_stream_act_local_4 <= conv2d_24_stream_act_local_4 + cparam_conv2d_24_inc_act_laddr_small;
          end 
          if((conv2d_24_col_select == 0)? cparam_conv2d_24_inc_act_laddr_conds_12 : 
          (conv2d_24_col_select == 1)? cparam_conv2d_24_inc_act_laddr_conds_13 : 
          (conv2d_24_col_select == 2)? cparam_conv2d_24_inc_act_laddr_conds_14 : 0) begin
            conv2d_24_stream_act_local_4 <= conv2d_24_stream_act_local_4 + cparam_conv2d_24_inc_act_laddr_large;
          end 
          if(conv2d_24_col_count >= cparam_conv2d_24_max_col_count) begin
            conv2d_24_stream_act_local_4 <= 0;
          end 
          if((conv2d_24_col_count >= cparam_conv2d_24_max_col_count) && cparam_conv2d_24_stream_act_local_small_flags_1) begin
            conv2d_24_stream_act_local_4 <= cparam_conv2d_24_stream_act_local_small_offset;
          end 
          if((conv2d_24_col_count >= cparam_conv2d_24_max_col_count) && cparam_conv2d_24_stream_act_local_large_flags_1) begin
            conv2d_24_stream_act_local_4 <= cparam_conv2d_24_stream_act_local_large_offset;
          end 
          if(!((conv2d_24_col_select == 0)? cparam_conv2d_24_inc_act_laddr_conds_15 : 
          (conv2d_24_col_select == 1)? cparam_conv2d_24_inc_act_laddr_conds_16 : 
          (conv2d_24_col_select == 2)? cparam_conv2d_24_inc_act_laddr_conds_17 : 0)) begin
            conv2d_24_stream_act_local_5 <= conv2d_24_stream_act_local_5 + cparam_conv2d_24_inc_act_laddr_small;
          end 
          if((conv2d_24_col_select == 0)? cparam_conv2d_24_inc_act_laddr_conds_15 : 
          (conv2d_24_col_select == 1)? cparam_conv2d_24_inc_act_laddr_conds_16 : 
          (conv2d_24_col_select == 2)? cparam_conv2d_24_inc_act_laddr_conds_17 : 0) begin
            conv2d_24_stream_act_local_5 <= conv2d_24_stream_act_local_5 + cparam_conv2d_24_inc_act_laddr_large;
          end 
          if(conv2d_24_col_count >= cparam_conv2d_24_max_col_count) begin
            conv2d_24_stream_act_local_5 <= 0;
          end 
          if((conv2d_24_col_count >= cparam_conv2d_24_max_col_count) && cparam_conv2d_24_stream_act_local_small_flags_2) begin
            conv2d_24_stream_act_local_5 <= cparam_conv2d_24_stream_act_local_small_offset;
          end 
          if((conv2d_24_col_count >= cparam_conv2d_24_max_col_count) && cparam_conv2d_24_stream_act_local_large_flags_2) begin
            conv2d_24_stream_act_local_5 <= cparam_conv2d_24_stream_act_local_large_offset;
          end 
          if(!((conv2d_24_col_select == 0)? cparam_conv2d_24_inc_act_laddr_conds_18 : 
          (conv2d_24_col_select == 1)? cparam_conv2d_24_inc_act_laddr_conds_19 : 
          (conv2d_24_col_select == 2)? cparam_conv2d_24_inc_act_laddr_conds_20 : 0)) begin
            conv2d_24_stream_act_local_6 <= conv2d_24_stream_act_local_6 + cparam_conv2d_24_inc_act_laddr_small;
          end 
          if((conv2d_24_col_select == 0)? cparam_conv2d_24_inc_act_laddr_conds_18 : 
          (conv2d_24_col_select == 1)? cparam_conv2d_24_inc_act_laddr_conds_19 : 
          (conv2d_24_col_select == 2)? cparam_conv2d_24_inc_act_laddr_conds_20 : 0) begin
            conv2d_24_stream_act_local_6 <= conv2d_24_stream_act_local_6 + cparam_conv2d_24_inc_act_laddr_large;
          end 
          if(conv2d_24_col_count >= cparam_conv2d_24_max_col_count) begin
            conv2d_24_stream_act_local_6 <= 0;
          end 
          if((conv2d_24_col_count >= cparam_conv2d_24_max_col_count) && cparam_conv2d_24_stream_act_local_small_flags_0) begin
            conv2d_24_stream_act_local_6 <= cparam_conv2d_24_stream_act_local_small_offset;
          end 
          if((conv2d_24_col_count >= cparam_conv2d_24_max_col_count) && cparam_conv2d_24_stream_act_local_large_flags_0) begin
            conv2d_24_stream_act_local_6 <= cparam_conv2d_24_stream_act_local_large_offset;
          end 
          if(!((conv2d_24_col_select == 0)? cparam_conv2d_24_inc_act_laddr_conds_21 : 
          (conv2d_24_col_select == 1)? cparam_conv2d_24_inc_act_laddr_conds_22 : 
          (conv2d_24_col_select == 2)? cparam_conv2d_24_inc_act_laddr_conds_23 : 0)) begin
            conv2d_24_stream_act_local_7 <= conv2d_24_stream_act_local_7 + cparam_conv2d_24_inc_act_laddr_small;
          end 
          if((conv2d_24_col_select == 0)? cparam_conv2d_24_inc_act_laddr_conds_21 : 
          (conv2d_24_col_select == 1)? cparam_conv2d_24_inc_act_laddr_conds_22 : 
          (conv2d_24_col_select == 2)? cparam_conv2d_24_inc_act_laddr_conds_23 : 0) begin
            conv2d_24_stream_act_local_7 <= conv2d_24_stream_act_local_7 + cparam_conv2d_24_inc_act_laddr_large;
          end 
          if(conv2d_24_col_count >= cparam_conv2d_24_max_col_count) begin
            conv2d_24_stream_act_local_7 <= 0;
          end 
          if((conv2d_24_col_count >= cparam_conv2d_24_max_col_count) && cparam_conv2d_24_stream_act_local_small_flags_1) begin
            conv2d_24_stream_act_local_7 <= cparam_conv2d_24_stream_act_local_small_offset;
          end 
          if((conv2d_24_col_count >= cparam_conv2d_24_max_col_count) && cparam_conv2d_24_stream_act_local_large_flags_1) begin
            conv2d_24_stream_act_local_7 <= cparam_conv2d_24_stream_act_local_large_offset;
          end 
          if(!((conv2d_24_col_select == 0)? cparam_conv2d_24_inc_act_laddr_conds_24 : 
          (conv2d_24_col_select == 1)? cparam_conv2d_24_inc_act_laddr_conds_25 : 
          (conv2d_24_col_select == 2)? cparam_conv2d_24_inc_act_laddr_conds_26 : 0)) begin
            conv2d_24_stream_act_local_8 <= conv2d_24_stream_act_local_8 + cparam_conv2d_24_inc_act_laddr_small;
          end 
          if((conv2d_24_col_select == 0)? cparam_conv2d_24_inc_act_laddr_conds_24 : 
          (conv2d_24_col_select == 1)? cparam_conv2d_24_inc_act_laddr_conds_25 : 
          (conv2d_24_col_select == 2)? cparam_conv2d_24_inc_act_laddr_conds_26 : 0) begin
            conv2d_24_stream_act_local_8 <= conv2d_24_stream_act_local_8 + cparam_conv2d_24_inc_act_laddr_large;
          end 
          if(conv2d_24_col_count >= cparam_conv2d_24_max_col_count) begin
            conv2d_24_stream_act_local_8 <= 0;
          end 
          if((conv2d_24_col_count >= cparam_conv2d_24_max_col_count) && cparam_conv2d_24_stream_act_local_small_flags_2) begin
            conv2d_24_stream_act_local_8 <= cparam_conv2d_24_stream_act_local_small_offset;
          end 
          if((conv2d_24_col_count >= cparam_conv2d_24_max_col_count) && cparam_conv2d_24_stream_act_local_large_flags_2) begin
            conv2d_24_stream_act_local_8 <= cparam_conv2d_24_stream_act_local_large_offset;
          end 
          if(cparam_conv2d_24_data_stationary == 0) begin
            conv2d_24_stream_out_local_col <= conv2d_24_stream_out_local_col + conv2d_24_next_stream_num_ops;
          end 
          if((cparam_conv2d_24_data_stationary == 0) && (conv2d_24_col_count >= cparam_conv2d_24_max_col_count)) begin
            conv2d_24_stream_out_local_col <= 0;
          end 
          if(cparam_conv2d_24_data_stationary == 1) begin
            conv2d_24_stream_out_local_col <= conv2d_24_stream_out_local_col + cparam_conv2d_24_inc_out_laddr_col;
          end 
          if((cparam_conv2d_24_data_stationary == 1) && (conv2d_24_col_count >= cparam_conv2d_24_max_col_count)) begin
            conv2d_24_stream_out_local_val <= conv2d_24_stream_out_local_val + conv2d_24_next_stream_num_ops;
            conv2d_24_stream_out_local_col <= 0;
          end 
          conv2d_24_col_count <= conv2d_24_col_count + cparam_conv2d_24_stride_col_par_col;
          if(conv2d_24_col_count >= cparam_conv2d_24_max_col_count) begin
            conv2d_24_col_count <= 0;
          end 
          conv2d_24_col_select <= conv2d_24_col_select + cparam_conv2d_24_stride_col_mod_filter_num;
          if(conv2d_24_col_select + cparam_conv2d_24_stride_col_mod_filter_num >= 3) begin
            conv2d_24_col_select <= conv2d_24_col_select - cparam_conv2d_24_filter_num_col_minus_stride_col_mod;
          end 
          if(conv2d_24_col_count >= cparam_conv2d_24_max_col_count) begin
            conv2d_24_col_select <= cparam_conv2d_24_col_select_initval;
          end 
          conv2d_24_comp_fsm <= conv2d_24_comp_fsm_2;
          if(conv2d_24_col_count >= cparam_conv2d_24_max_col_count) begin
            conv2d_24_comp_fsm <= conv2d_24_comp_fsm_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_24_source_7_source_pat_fsm_0_1 = 1;
  localparam _stream_conv2d_24_source_7_source_pat_fsm_0_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_24_source_7_source_pat_fsm_0 <= _stream_conv2d_24_source_7_source_pat_fsm_0_init;
    end else begin
      case(_stream_conv2d_24_source_7_source_pat_fsm_0)
        _stream_conv2d_24_source_7_source_pat_fsm_0_init: begin
          if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_7_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_7_source_pat_fsm_0 <= _stream_conv2d_24_source_7_source_pat_fsm_0_1;
          end 
        end
        _stream_conv2d_24_source_7_source_pat_fsm_0_1: begin
          if(_stream_conv2d_24_source_stop && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_7_source_pat_fsm_0 <= _stream_conv2d_24_source_7_source_pat_fsm_0_init;
          end 
          if((_source_stream_conv2d_24_source_7_pat_count_0 == 0) && (_source_stream_conv2d_24_source_7_pat_count_1 == 0) && (_source_stream_conv2d_24_source_7_pat_count_2 == 0) && (_source_stream_conv2d_24_source_7_pat_count_3 == 0) && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_7_source_pat_fsm_0 <= _stream_conv2d_24_source_7_source_pat_fsm_0_2;
          end 
        end
        _stream_conv2d_24_source_7_source_pat_fsm_0_2: begin
          if(_stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_7_source_pat_fsm_0 <= _stream_conv2d_24_source_7_source_pat_fsm_0_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_409 <= 0;
      _tmp_1668 <= 0;
    end else begin
      if(_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_9_source_ram_renable && (_stream_conv2d_24_source_9_source_sel == 2)) begin
        _tmp_409 <= read_rtl_bank_408;
      end 
      if(_stream_matmul_55_stream_oready && _stream_matmul_55_source_9_source_ram_renable && (_stream_matmul_55_source_9_source_sel == 2)) begin
        _tmp_1668 <= read_rtl_bank_1667;
      end 
    end
  end

  localparam _stream_conv2d_24_source_9_source_pat_fsm_1_1 = 1;
  localparam _stream_conv2d_24_source_9_source_pat_fsm_1_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_24_source_9_source_pat_fsm_1 <= _stream_conv2d_24_source_9_source_pat_fsm_1_init;
    end else begin
      case(_stream_conv2d_24_source_9_source_pat_fsm_1)
        _stream_conv2d_24_source_9_source_pat_fsm_1_init: begin
          if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_9_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_9_source_pat_fsm_1 <= _stream_conv2d_24_source_9_source_pat_fsm_1_1;
          end 
        end
        _stream_conv2d_24_source_9_source_pat_fsm_1_1: begin
          if(_stream_conv2d_24_source_stop && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_9_source_pat_fsm_1 <= _stream_conv2d_24_source_9_source_pat_fsm_1_init;
          end 
          if((_source_stream_conv2d_24_source_9_pat_count_0 == 0) && (_source_stream_conv2d_24_source_9_pat_count_1 == 0) && (_source_stream_conv2d_24_source_9_pat_count_2 == 0) && (_source_stream_conv2d_24_source_9_pat_count_3 == 0) && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_9_source_pat_fsm_1 <= _stream_conv2d_24_source_9_source_pat_fsm_1_2;
          end 
        end
        _stream_conv2d_24_source_9_source_pat_fsm_1_2: begin
          if(_stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_9_source_pat_fsm_1 <= _stream_conv2d_24_source_9_source_pat_fsm_1_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_432 <= 0;
      _tmp_1496 <= 0;
    end else begin
      if(_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_20_source_ram_renable && (_stream_conv2d_24_source_20_source_sel == 3)) begin
        _tmp_432 <= read_rtl_bank_431;
      end 
      if(_stream_avg_pool_serial_52_stream_oready && _stream_avg_pool_serial_52_source_1_source_ram_renable && (_stream_avg_pool_serial_52_source_1_source_sel == 1)) begin
        _tmp_1496 <= read_rtl_bank_1495;
      end 
    end
  end

  localparam _stream_conv2d_24_source_20_source_pat_fsm_2_1 = 1;
  localparam _stream_conv2d_24_source_20_source_pat_fsm_2_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_24_source_20_source_pat_fsm_2 <= _stream_conv2d_24_source_20_source_pat_fsm_2_init;
    end else begin
      case(_stream_conv2d_24_source_20_source_pat_fsm_2)
        _stream_conv2d_24_source_20_source_pat_fsm_2_init: begin
          if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_20_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_20_source_pat_fsm_2 <= _stream_conv2d_24_source_20_source_pat_fsm_2_1;
          end 
        end
        _stream_conv2d_24_source_20_source_pat_fsm_2_1: begin
          if(_stream_conv2d_24_source_stop && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_20_source_pat_fsm_2 <= _stream_conv2d_24_source_20_source_pat_fsm_2_init;
          end 
          if((_source_stream_conv2d_24_source_20_pat_count_0 == 0) && (_source_stream_conv2d_24_source_20_pat_count_1 == 0) && (_source_stream_conv2d_24_source_20_pat_count_2 == 0) && (_source_stream_conv2d_24_source_20_pat_count_3 == 0) && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_20_source_pat_fsm_2 <= _stream_conv2d_24_source_20_source_pat_fsm_2_2;
          end 
        end
        _stream_conv2d_24_source_20_source_pat_fsm_2_2: begin
          if(_stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_20_source_pat_fsm_2 <= _stream_conv2d_24_source_20_source_pat_fsm_2_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_445 <= 0;
    end else begin
      if(_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_21_source_ram_renable && (_stream_conv2d_24_source_21_source_sel == 4)) begin
        _tmp_445 <= read_rtl_bank_444;
      end 
    end
  end

  localparam _stream_conv2d_24_source_21_source_pat_fsm_3_1 = 1;
  localparam _stream_conv2d_24_source_21_source_pat_fsm_3_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_24_source_21_source_pat_fsm_3 <= _stream_conv2d_24_source_21_source_pat_fsm_3_init;
    end else begin
      case(_stream_conv2d_24_source_21_source_pat_fsm_3)
        _stream_conv2d_24_source_21_source_pat_fsm_3_init: begin
          if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_21_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_21_source_pat_fsm_3 <= _stream_conv2d_24_source_21_source_pat_fsm_3_1;
          end 
        end
        _stream_conv2d_24_source_21_source_pat_fsm_3_1: begin
          if(_stream_conv2d_24_source_stop && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_21_source_pat_fsm_3 <= _stream_conv2d_24_source_21_source_pat_fsm_3_init;
          end 
          if((_source_stream_conv2d_24_source_21_pat_count_0 == 0) && (_source_stream_conv2d_24_source_21_pat_count_1 == 0) && (_source_stream_conv2d_24_source_21_pat_count_2 == 0) && (_source_stream_conv2d_24_source_21_pat_count_3 == 0) && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_21_source_pat_fsm_3 <= _stream_conv2d_24_source_21_source_pat_fsm_3_2;
          end 
        end
        _stream_conv2d_24_source_21_source_pat_fsm_3_2: begin
          if(_stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_21_source_pat_fsm_3 <= _stream_conv2d_24_source_21_source_pat_fsm_3_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_458 <= 0;
    end else begin
      if(_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_22_source_ram_renable && (_stream_conv2d_24_source_22_source_sel == 5)) begin
        _tmp_458 <= read_rtl_bank_457;
      end 
    end
  end

  localparam _stream_conv2d_24_source_22_source_pat_fsm_4_1 = 1;
  localparam _stream_conv2d_24_source_22_source_pat_fsm_4_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_24_source_22_source_pat_fsm_4 <= _stream_conv2d_24_source_22_source_pat_fsm_4_init;
    end else begin
      case(_stream_conv2d_24_source_22_source_pat_fsm_4)
        _stream_conv2d_24_source_22_source_pat_fsm_4_init: begin
          if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_22_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_22_source_pat_fsm_4 <= _stream_conv2d_24_source_22_source_pat_fsm_4_1;
          end 
        end
        _stream_conv2d_24_source_22_source_pat_fsm_4_1: begin
          if(_stream_conv2d_24_source_stop && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_22_source_pat_fsm_4 <= _stream_conv2d_24_source_22_source_pat_fsm_4_init;
          end 
          if((_source_stream_conv2d_24_source_22_pat_count_0 == 0) && (_source_stream_conv2d_24_source_22_pat_count_1 == 0) && (_source_stream_conv2d_24_source_22_pat_count_2 == 0) && (_source_stream_conv2d_24_source_22_pat_count_3 == 0) && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_22_source_pat_fsm_4 <= _stream_conv2d_24_source_22_source_pat_fsm_4_2;
          end 
        end
        _stream_conv2d_24_source_22_source_pat_fsm_4_2: begin
          if(_stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_22_source_pat_fsm_4 <= _stream_conv2d_24_source_22_source_pat_fsm_4_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_471 <= 0;
    end else begin
      if(_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_23_source_ram_renable && (_stream_conv2d_24_source_23_source_sel == 6)) begin
        _tmp_471 <= read_rtl_bank_470;
      end 
    end
  end

  localparam _stream_conv2d_24_source_23_source_pat_fsm_5_1 = 1;
  localparam _stream_conv2d_24_source_23_source_pat_fsm_5_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_24_source_23_source_pat_fsm_5 <= _stream_conv2d_24_source_23_source_pat_fsm_5_init;
    end else begin
      case(_stream_conv2d_24_source_23_source_pat_fsm_5)
        _stream_conv2d_24_source_23_source_pat_fsm_5_init: begin
          if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_23_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_23_source_pat_fsm_5 <= _stream_conv2d_24_source_23_source_pat_fsm_5_1;
          end 
        end
        _stream_conv2d_24_source_23_source_pat_fsm_5_1: begin
          if(_stream_conv2d_24_source_stop && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_23_source_pat_fsm_5 <= _stream_conv2d_24_source_23_source_pat_fsm_5_init;
          end 
          if((_source_stream_conv2d_24_source_23_pat_count_0 == 0) && (_source_stream_conv2d_24_source_23_pat_count_1 == 0) && (_source_stream_conv2d_24_source_23_pat_count_2 == 0) && (_source_stream_conv2d_24_source_23_pat_count_3 == 0) && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_23_source_pat_fsm_5 <= _stream_conv2d_24_source_23_source_pat_fsm_5_2;
          end 
        end
        _stream_conv2d_24_source_23_source_pat_fsm_5_2: begin
          if(_stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_23_source_pat_fsm_5 <= _stream_conv2d_24_source_23_source_pat_fsm_5_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_484 <= 0;
    end else begin
      if(_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_24_source_ram_renable && (_stream_conv2d_24_source_24_source_sel == 7)) begin
        _tmp_484 <= read_rtl_bank_483;
      end 
    end
  end

  localparam _stream_conv2d_24_source_24_source_pat_fsm_6_1 = 1;
  localparam _stream_conv2d_24_source_24_source_pat_fsm_6_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_24_source_24_source_pat_fsm_6 <= _stream_conv2d_24_source_24_source_pat_fsm_6_init;
    end else begin
      case(_stream_conv2d_24_source_24_source_pat_fsm_6)
        _stream_conv2d_24_source_24_source_pat_fsm_6_init: begin
          if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_24_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_24_source_pat_fsm_6 <= _stream_conv2d_24_source_24_source_pat_fsm_6_1;
          end 
        end
        _stream_conv2d_24_source_24_source_pat_fsm_6_1: begin
          if(_stream_conv2d_24_source_stop && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_24_source_pat_fsm_6 <= _stream_conv2d_24_source_24_source_pat_fsm_6_init;
          end 
          if((_source_stream_conv2d_24_source_24_pat_count_0 == 0) && (_source_stream_conv2d_24_source_24_pat_count_1 == 0) && (_source_stream_conv2d_24_source_24_pat_count_2 == 0) && (_source_stream_conv2d_24_source_24_pat_count_3 == 0) && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_24_source_pat_fsm_6 <= _stream_conv2d_24_source_24_source_pat_fsm_6_2;
          end 
        end
        _stream_conv2d_24_source_24_source_pat_fsm_6_2: begin
          if(_stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_24_source_pat_fsm_6 <= _stream_conv2d_24_source_24_source_pat_fsm_6_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_497 <= 0;
    end else begin
      if(_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_25_source_ram_renable && (_stream_conv2d_24_source_25_source_sel == 8)) begin
        _tmp_497 <= read_rtl_bank_496;
      end 
    end
  end

  localparam _stream_conv2d_24_source_25_source_pat_fsm_7_1 = 1;
  localparam _stream_conv2d_24_source_25_source_pat_fsm_7_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_24_source_25_source_pat_fsm_7 <= _stream_conv2d_24_source_25_source_pat_fsm_7_init;
    end else begin
      case(_stream_conv2d_24_source_25_source_pat_fsm_7)
        _stream_conv2d_24_source_25_source_pat_fsm_7_init: begin
          if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_25_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_25_source_pat_fsm_7 <= _stream_conv2d_24_source_25_source_pat_fsm_7_1;
          end 
        end
        _stream_conv2d_24_source_25_source_pat_fsm_7_1: begin
          if(_stream_conv2d_24_source_stop && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_25_source_pat_fsm_7 <= _stream_conv2d_24_source_25_source_pat_fsm_7_init;
          end 
          if((_source_stream_conv2d_24_source_25_pat_count_0 == 0) && (_source_stream_conv2d_24_source_25_pat_count_1 == 0) && (_source_stream_conv2d_24_source_25_pat_count_2 == 0) && (_source_stream_conv2d_24_source_25_pat_count_3 == 0) && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_25_source_pat_fsm_7 <= _stream_conv2d_24_source_25_source_pat_fsm_7_2;
          end 
        end
        _stream_conv2d_24_source_25_source_pat_fsm_7_2: begin
          if(_stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_25_source_pat_fsm_7 <= _stream_conv2d_24_source_25_source_pat_fsm_7_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_510 <= 0;
    end else begin
      if(_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_26_source_ram_renable && (_stream_conv2d_24_source_26_source_sel == 9)) begin
        _tmp_510 <= read_rtl_bank_509;
      end 
    end
  end

  localparam _stream_conv2d_24_source_26_source_pat_fsm_8_1 = 1;
  localparam _stream_conv2d_24_source_26_source_pat_fsm_8_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_24_source_26_source_pat_fsm_8 <= _stream_conv2d_24_source_26_source_pat_fsm_8_init;
    end else begin
      case(_stream_conv2d_24_source_26_source_pat_fsm_8)
        _stream_conv2d_24_source_26_source_pat_fsm_8_init: begin
          if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_26_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_26_source_pat_fsm_8 <= _stream_conv2d_24_source_26_source_pat_fsm_8_1;
          end 
        end
        _stream_conv2d_24_source_26_source_pat_fsm_8_1: begin
          if(_stream_conv2d_24_source_stop && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_26_source_pat_fsm_8 <= _stream_conv2d_24_source_26_source_pat_fsm_8_init;
          end 
          if((_source_stream_conv2d_24_source_26_pat_count_0 == 0) && (_source_stream_conv2d_24_source_26_pat_count_1 == 0) && (_source_stream_conv2d_24_source_26_pat_count_2 == 0) && (_source_stream_conv2d_24_source_26_pat_count_3 == 0) && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_26_source_pat_fsm_8 <= _stream_conv2d_24_source_26_source_pat_fsm_8_2;
          end 
        end
        _stream_conv2d_24_source_26_source_pat_fsm_8_2: begin
          if(_stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_26_source_pat_fsm_8 <= _stream_conv2d_24_source_26_source_pat_fsm_8_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_523 <= 0;
    end else begin
      if(_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_27_source_ram_renable && (_stream_conv2d_24_source_27_source_sel == 10)) begin
        _tmp_523 <= read_rtl_bank_522;
      end 
    end
  end

  localparam _stream_conv2d_24_source_27_source_pat_fsm_9_1 = 1;
  localparam _stream_conv2d_24_source_27_source_pat_fsm_9_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_24_source_27_source_pat_fsm_9 <= _stream_conv2d_24_source_27_source_pat_fsm_9_init;
    end else begin
      case(_stream_conv2d_24_source_27_source_pat_fsm_9)
        _stream_conv2d_24_source_27_source_pat_fsm_9_init: begin
          if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_27_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_27_source_pat_fsm_9 <= _stream_conv2d_24_source_27_source_pat_fsm_9_1;
          end 
        end
        _stream_conv2d_24_source_27_source_pat_fsm_9_1: begin
          if(_stream_conv2d_24_source_stop && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_27_source_pat_fsm_9 <= _stream_conv2d_24_source_27_source_pat_fsm_9_init;
          end 
          if((_source_stream_conv2d_24_source_27_pat_count_0 == 0) && (_source_stream_conv2d_24_source_27_pat_count_1 == 0) && (_source_stream_conv2d_24_source_27_pat_count_2 == 0) && (_source_stream_conv2d_24_source_27_pat_count_3 == 0) && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_27_source_pat_fsm_9 <= _stream_conv2d_24_source_27_source_pat_fsm_9_2;
          end 
        end
        _stream_conv2d_24_source_27_source_pat_fsm_9_2: begin
          if(_stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_27_source_pat_fsm_9 <= _stream_conv2d_24_source_27_source_pat_fsm_9_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_536 <= 0;
    end else begin
      if(_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_28_source_ram_renable && (_stream_conv2d_24_source_28_source_sel == 11)) begin
        _tmp_536 <= read_rtl_bank_535;
      end 
    end
  end

  localparam _stream_conv2d_24_source_28_source_pat_fsm_10_1 = 1;
  localparam _stream_conv2d_24_source_28_source_pat_fsm_10_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_24_source_28_source_pat_fsm_10 <= _stream_conv2d_24_source_28_source_pat_fsm_10_init;
    end else begin
      case(_stream_conv2d_24_source_28_source_pat_fsm_10)
        _stream_conv2d_24_source_28_source_pat_fsm_10_init: begin
          if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_28_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_28_source_pat_fsm_10 <= _stream_conv2d_24_source_28_source_pat_fsm_10_1;
          end 
        end
        _stream_conv2d_24_source_28_source_pat_fsm_10_1: begin
          if(_stream_conv2d_24_source_stop && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_28_source_pat_fsm_10 <= _stream_conv2d_24_source_28_source_pat_fsm_10_init;
          end 
          if((_source_stream_conv2d_24_source_28_pat_count_0 == 0) && (_source_stream_conv2d_24_source_28_pat_count_1 == 0) && (_source_stream_conv2d_24_source_28_pat_count_2 == 0) && (_source_stream_conv2d_24_source_28_pat_count_3 == 0) && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_28_source_pat_fsm_10 <= _stream_conv2d_24_source_28_source_pat_fsm_10_2;
          end 
        end
        _stream_conv2d_24_source_28_source_pat_fsm_10_2: begin
          if(_stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_28_source_pat_fsm_10 <= _stream_conv2d_24_source_28_source_pat_fsm_10_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_549 <= 0;
    end else begin
      if(_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_29_source_ram_renable && (_stream_conv2d_24_source_29_source_sel == 12)) begin
        _tmp_549 <= read_rtl_bank_548;
      end 
    end
  end

  localparam _stream_conv2d_24_source_29_source_pat_fsm_11_1 = 1;
  localparam _stream_conv2d_24_source_29_source_pat_fsm_11_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_24_source_29_source_pat_fsm_11 <= _stream_conv2d_24_source_29_source_pat_fsm_11_init;
    end else begin
      case(_stream_conv2d_24_source_29_source_pat_fsm_11)
        _stream_conv2d_24_source_29_source_pat_fsm_11_init: begin
          if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_29_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_29_source_pat_fsm_11 <= _stream_conv2d_24_source_29_source_pat_fsm_11_1;
          end 
        end
        _stream_conv2d_24_source_29_source_pat_fsm_11_1: begin
          if(_stream_conv2d_24_source_stop && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_29_source_pat_fsm_11 <= _stream_conv2d_24_source_29_source_pat_fsm_11_init;
          end 
          if((_source_stream_conv2d_24_source_29_pat_count_0 == 0) && (_source_stream_conv2d_24_source_29_pat_count_1 == 0) && (_source_stream_conv2d_24_source_29_pat_count_2 == 0) && (_source_stream_conv2d_24_source_29_pat_count_3 == 0) && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_29_source_pat_fsm_11 <= _stream_conv2d_24_source_29_source_pat_fsm_11_2;
          end 
        end
        _stream_conv2d_24_source_29_source_pat_fsm_11_2: begin
          if(_stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_29_source_pat_fsm_11 <= _stream_conv2d_24_source_29_source_pat_fsm_11_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_562 <= 0;
    end else begin
      if(_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_30_source_ram_renable && (_stream_conv2d_24_source_30_source_sel == 13)) begin
        _tmp_562 <= read_rtl_bank_561;
      end 
    end
  end

  localparam _stream_conv2d_24_source_30_source_pat_fsm_12_1 = 1;
  localparam _stream_conv2d_24_source_30_source_pat_fsm_12_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_24_source_30_source_pat_fsm_12 <= _stream_conv2d_24_source_30_source_pat_fsm_12_init;
    end else begin
      case(_stream_conv2d_24_source_30_source_pat_fsm_12)
        _stream_conv2d_24_source_30_source_pat_fsm_12_init: begin
          if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_30_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_30_source_pat_fsm_12 <= _stream_conv2d_24_source_30_source_pat_fsm_12_1;
          end 
        end
        _stream_conv2d_24_source_30_source_pat_fsm_12_1: begin
          if(_stream_conv2d_24_source_stop && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_30_source_pat_fsm_12 <= _stream_conv2d_24_source_30_source_pat_fsm_12_init;
          end 
          if((_source_stream_conv2d_24_source_30_pat_count_0 == 0) && (_source_stream_conv2d_24_source_30_pat_count_1 == 0) && (_source_stream_conv2d_24_source_30_pat_count_2 == 0) && (_source_stream_conv2d_24_source_30_pat_count_3 == 0) && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_30_source_pat_fsm_12 <= _stream_conv2d_24_source_30_source_pat_fsm_12_2;
          end 
        end
        _stream_conv2d_24_source_30_source_pat_fsm_12_2: begin
          if(_stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_30_source_pat_fsm_12 <= _stream_conv2d_24_source_30_source_pat_fsm_12_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_575 <= 0;
    end else begin
      if(_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_31_source_ram_renable && (_stream_conv2d_24_source_31_source_sel == 14)) begin
        _tmp_575 <= read_rtl_bank_574;
      end 
    end
  end

  localparam _stream_conv2d_24_source_31_source_pat_fsm_13_1 = 1;
  localparam _stream_conv2d_24_source_31_source_pat_fsm_13_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_24_source_31_source_pat_fsm_13 <= _stream_conv2d_24_source_31_source_pat_fsm_13_init;
    end else begin
      case(_stream_conv2d_24_source_31_source_pat_fsm_13)
        _stream_conv2d_24_source_31_source_pat_fsm_13_init: begin
          if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_31_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_31_source_pat_fsm_13 <= _stream_conv2d_24_source_31_source_pat_fsm_13_1;
          end 
        end
        _stream_conv2d_24_source_31_source_pat_fsm_13_1: begin
          if(_stream_conv2d_24_source_stop && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_31_source_pat_fsm_13 <= _stream_conv2d_24_source_31_source_pat_fsm_13_init;
          end 
          if((_source_stream_conv2d_24_source_31_pat_count_0 == 0) && (_source_stream_conv2d_24_source_31_pat_count_1 == 0) && (_source_stream_conv2d_24_source_31_pat_count_2 == 0) && (_source_stream_conv2d_24_source_31_pat_count_3 == 0) && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_31_source_pat_fsm_13 <= _stream_conv2d_24_source_31_source_pat_fsm_13_2;
          end 
        end
        _stream_conv2d_24_source_31_source_pat_fsm_13_2: begin
          if(_stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_31_source_pat_fsm_13 <= _stream_conv2d_24_source_31_source_pat_fsm_13_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_588 <= 0;
    end else begin
      if(_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_32_source_ram_renable && (_stream_conv2d_24_source_32_source_sel == 15)) begin
        _tmp_588 <= read_rtl_bank_587;
      end 
    end
  end

  localparam _stream_conv2d_24_source_32_source_pat_fsm_14_1 = 1;
  localparam _stream_conv2d_24_source_32_source_pat_fsm_14_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_24_source_32_source_pat_fsm_14 <= _stream_conv2d_24_source_32_source_pat_fsm_14_init;
    end else begin
      case(_stream_conv2d_24_source_32_source_pat_fsm_14)
        _stream_conv2d_24_source_32_source_pat_fsm_14_init: begin
          if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_32_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_32_source_pat_fsm_14 <= _stream_conv2d_24_source_32_source_pat_fsm_14_1;
          end 
        end
        _stream_conv2d_24_source_32_source_pat_fsm_14_1: begin
          if(_stream_conv2d_24_source_stop && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_32_source_pat_fsm_14 <= _stream_conv2d_24_source_32_source_pat_fsm_14_init;
          end 
          if((_source_stream_conv2d_24_source_32_pat_count_0 == 0) && (_source_stream_conv2d_24_source_32_pat_count_1 == 0) && (_source_stream_conv2d_24_source_32_pat_count_2 == 0) && (_source_stream_conv2d_24_source_32_pat_count_3 == 0) && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_32_source_pat_fsm_14 <= _stream_conv2d_24_source_32_source_pat_fsm_14_2;
          end 
        end
        _stream_conv2d_24_source_32_source_pat_fsm_14_2: begin
          if(_stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_32_source_pat_fsm_14 <= _stream_conv2d_24_source_32_source_pat_fsm_14_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_601 <= 0;
    end else begin
      if(_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_33_source_ram_renable && (_stream_conv2d_24_source_33_source_sel == 16)) begin
        _tmp_601 <= read_rtl_bank_600;
      end 
    end
  end

  localparam _stream_conv2d_24_source_33_source_pat_fsm_15_1 = 1;
  localparam _stream_conv2d_24_source_33_source_pat_fsm_15_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_24_source_33_source_pat_fsm_15 <= _stream_conv2d_24_source_33_source_pat_fsm_15_init;
    end else begin
      case(_stream_conv2d_24_source_33_source_pat_fsm_15)
        _stream_conv2d_24_source_33_source_pat_fsm_15_init: begin
          if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_33_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_33_source_pat_fsm_15 <= _stream_conv2d_24_source_33_source_pat_fsm_15_1;
          end 
        end
        _stream_conv2d_24_source_33_source_pat_fsm_15_1: begin
          if(_stream_conv2d_24_source_stop && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_33_source_pat_fsm_15 <= _stream_conv2d_24_source_33_source_pat_fsm_15_init;
          end 
          if((_source_stream_conv2d_24_source_33_pat_count_0 == 0) && (_source_stream_conv2d_24_source_33_pat_count_1 == 0) && (_source_stream_conv2d_24_source_33_pat_count_2 == 0) && (_source_stream_conv2d_24_source_33_pat_count_3 == 0) && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_33_source_pat_fsm_15 <= _stream_conv2d_24_source_33_source_pat_fsm_15_2;
          end 
        end
        _stream_conv2d_24_source_33_source_pat_fsm_15_2: begin
          if(_stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_33_source_pat_fsm_15 <= _stream_conv2d_24_source_33_source_pat_fsm_15_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_614 <= 0;
    end else begin
      if(_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_34_source_ram_renable && (_stream_conv2d_24_source_34_source_sel == 17)) begin
        _tmp_614 <= read_rtl_bank_613;
      end 
    end
  end

  localparam _stream_conv2d_24_source_34_source_pat_fsm_16_1 = 1;
  localparam _stream_conv2d_24_source_34_source_pat_fsm_16_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_24_source_34_source_pat_fsm_16 <= _stream_conv2d_24_source_34_source_pat_fsm_16_init;
    end else begin
      case(_stream_conv2d_24_source_34_source_pat_fsm_16)
        _stream_conv2d_24_source_34_source_pat_fsm_16_init: begin
          if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_34_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_34_source_pat_fsm_16 <= _stream_conv2d_24_source_34_source_pat_fsm_16_1;
          end 
        end
        _stream_conv2d_24_source_34_source_pat_fsm_16_1: begin
          if(_stream_conv2d_24_source_stop && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_34_source_pat_fsm_16 <= _stream_conv2d_24_source_34_source_pat_fsm_16_init;
          end 
          if((_source_stream_conv2d_24_source_34_pat_count_0 == 0) && (_source_stream_conv2d_24_source_34_pat_count_1 == 0) && (_source_stream_conv2d_24_source_34_pat_count_2 == 0) && (_source_stream_conv2d_24_source_34_pat_count_3 == 0) && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_34_source_pat_fsm_16 <= _stream_conv2d_24_source_34_source_pat_fsm_16_2;
          end 
        end
        _stream_conv2d_24_source_34_source_pat_fsm_16_2: begin
          if(_stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_34_source_pat_fsm_16 <= _stream_conv2d_24_source_34_source_pat_fsm_16_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_627 <= 0;
    end else begin
      if(_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_35_source_ram_renable && (_stream_conv2d_24_source_35_source_sel == 18)) begin
        _tmp_627 <= read_rtl_bank_626;
      end 
    end
  end

  localparam _stream_conv2d_24_source_35_source_pat_fsm_17_1 = 1;
  localparam _stream_conv2d_24_source_35_source_pat_fsm_17_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_24_source_35_source_pat_fsm_17 <= _stream_conv2d_24_source_35_source_pat_fsm_17_init;
    end else begin
      case(_stream_conv2d_24_source_35_source_pat_fsm_17)
        _stream_conv2d_24_source_35_source_pat_fsm_17_init: begin
          if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_35_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_35_source_pat_fsm_17 <= _stream_conv2d_24_source_35_source_pat_fsm_17_1;
          end 
        end
        _stream_conv2d_24_source_35_source_pat_fsm_17_1: begin
          if(_stream_conv2d_24_source_stop && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_35_source_pat_fsm_17 <= _stream_conv2d_24_source_35_source_pat_fsm_17_init;
          end 
          if((_source_stream_conv2d_24_source_35_pat_count_0 == 0) && (_source_stream_conv2d_24_source_35_pat_count_1 == 0) && (_source_stream_conv2d_24_source_35_pat_count_2 == 0) && (_source_stream_conv2d_24_source_35_pat_count_3 == 0) && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_35_source_pat_fsm_17 <= _stream_conv2d_24_source_35_source_pat_fsm_17_2;
          end 
        end
        _stream_conv2d_24_source_35_source_pat_fsm_17_2: begin
          if(_stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_35_source_pat_fsm_17 <= _stream_conv2d_24_source_35_source_pat_fsm_17_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_640 <= 0;
    end else begin
      if(_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_36_source_ram_renable && (_stream_conv2d_24_source_36_source_sel == 19)) begin
        _tmp_640 <= read_rtl_bank_639;
      end 
    end
  end

  localparam _stream_conv2d_24_source_36_source_pat_fsm_18_1 = 1;
  localparam _stream_conv2d_24_source_36_source_pat_fsm_18_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_24_source_36_source_pat_fsm_18 <= _stream_conv2d_24_source_36_source_pat_fsm_18_init;
    end else begin
      case(_stream_conv2d_24_source_36_source_pat_fsm_18)
        _stream_conv2d_24_source_36_source_pat_fsm_18_init: begin
          if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_36_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_36_source_pat_fsm_18 <= _stream_conv2d_24_source_36_source_pat_fsm_18_1;
          end 
        end
        _stream_conv2d_24_source_36_source_pat_fsm_18_1: begin
          if(_stream_conv2d_24_source_stop && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_36_source_pat_fsm_18 <= _stream_conv2d_24_source_36_source_pat_fsm_18_init;
          end 
          if((_source_stream_conv2d_24_source_36_pat_count_0 == 0) && (_source_stream_conv2d_24_source_36_pat_count_1 == 0) && (_source_stream_conv2d_24_source_36_pat_count_2 == 0) && (_source_stream_conv2d_24_source_36_pat_count_3 == 0) && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_36_source_pat_fsm_18 <= _stream_conv2d_24_source_36_source_pat_fsm_18_2;
          end 
        end
        _stream_conv2d_24_source_36_source_pat_fsm_18_2: begin
          if(_stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_36_source_pat_fsm_18 <= _stream_conv2d_24_source_36_source_pat_fsm_18_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_653 <= 0;
    end else begin
      if(_stream_conv2d_24_stream_oready && _stream_conv2d_24_source_37_source_ram_renable && (_stream_conv2d_24_source_37_source_sel == 20)) begin
        _tmp_653 <= read_rtl_bank_652;
      end 
    end
  end

  localparam _stream_conv2d_24_source_37_source_pat_fsm_19_1 = 1;
  localparam _stream_conv2d_24_source_37_source_pat_fsm_19_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_24_source_37_source_pat_fsm_19 <= _stream_conv2d_24_source_37_source_pat_fsm_19_init;
    end else begin
      case(_stream_conv2d_24_source_37_source_pat_fsm_19)
        _stream_conv2d_24_source_37_source_pat_fsm_19_init: begin
          if(_stream_conv2d_24_source_start && _stream_conv2d_24_source_37_source_mode & 5'b10 && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_37_source_pat_fsm_19 <= _stream_conv2d_24_source_37_source_pat_fsm_19_1;
          end 
        end
        _stream_conv2d_24_source_37_source_pat_fsm_19_1: begin
          if(_stream_conv2d_24_source_stop && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_37_source_pat_fsm_19 <= _stream_conv2d_24_source_37_source_pat_fsm_19_init;
          end 
          if((_source_stream_conv2d_24_source_37_pat_count_0 == 0) && (_source_stream_conv2d_24_source_37_pat_count_1 == 0) && (_source_stream_conv2d_24_source_37_pat_count_2 == 0) && (_source_stream_conv2d_24_source_37_pat_count_3 == 0) && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_37_source_pat_fsm_19 <= _stream_conv2d_24_source_37_source_pat_fsm_19_2;
          end 
        end
        _stream_conv2d_24_source_37_source_pat_fsm_19_2: begin
          if(_stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_source_37_source_pat_fsm_19 <= _stream_conv2d_24_source_37_source_pat_fsm_19_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_24_sink_50_sink_fsm_20_1 = 1;
  localparam _stream_conv2d_24_sink_50_sink_fsm_20_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_24_sink_50_sink_fsm_20 <= _stream_conv2d_24_sink_50_sink_fsm_20_init;
    end else begin
      case(_stream_conv2d_24_sink_50_sink_fsm_20)
        _stream_conv2d_24_sink_50_sink_fsm_20_init: begin
          if(_stream_conv2d_24_sink_start && _stream_conv2d_24_sink_50_sink_mode & 5'b1 && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_sink_50_sink_fsm_20 <= _stream_conv2d_24_sink_50_sink_fsm_20_1;
          end 
        end
        _stream_conv2d_24_sink_50_sink_fsm_20_1: begin
          if(_stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_sink_50_sink_fsm_20 <= _stream_conv2d_24_sink_50_sink_fsm_20_2;
          end 
        end
        _stream_conv2d_24_sink_50_sink_fsm_20_2: begin
          if(stream_conv2d_24_sink_51_data && (_stream_conv2d_24_sink_50_sink_count == 1) && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_sink_50_sink_fsm_20 <= _stream_conv2d_24_sink_50_sink_fsm_20_init;
          end 
          if(_stream_conv2d_24_sink_stop && _stream_conv2d_24_stream_oready) begin
            _stream_conv2d_24_sink_50_sink_fsm_20 <= _stream_conv2d_24_sink_50_sink_fsm_20_init;
          end 
        end
      endcase
    end
  end

  localparam _maxi_write_req_fsm_1 = 1;

  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      _maxi_write_req_fsm <= _maxi_write_req_fsm_init;
      _maxi_write_cont <= 0;
    end else begin
      case(_maxi_write_req_fsm)
        _maxi_write_req_fsm_init: begin
          if((_maxi_write_req_fsm == 0) && (_maxi_write_start || _maxi_write_cont) && !_maxi_write_req_fifo_almost_full) begin
            _maxi_write_req_fsm <= _maxi_write_req_fsm_1;
          end 
        end
        _maxi_write_req_fsm_1: begin
          if((_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (maxi_awready || !maxi_awvalid) && (_maxi_outstanding_wcount < 6)) begin
            _maxi_write_cont <= 1;
          end 
          if((_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (maxi_awready || !maxi_awvalid) && (_maxi_outstanding_wcount < 6) && (_maxi_write_global_size == 0)) begin
            _maxi_write_cont <= 0;
          end 
          if((_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (maxi_awready || !maxi_awvalid) && (_maxi_outstanding_wcount < 6)) begin
            _maxi_write_req_fsm <= _maxi_write_req_fsm_init;
          end 
        end
      endcase
    end
  end

  localparam _maxi_write_data_fsm_1 = 1;
  localparam _maxi_write_data_fsm_2 = 2;

  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      _maxi_write_data_fsm <= _maxi_write_data_fsm_init;
    end else begin
      case(_maxi_write_data_fsm)
        _maxi_write_data_fsm_init: begin
          if(!_maxi_write_data_busy && !_maxi_write_req_fifo_empty && (_maxi_write_op_sel_fifo == 1)) begin
            _maxi_write_data_fsm <= _maxi_write_data_fsm_1;
          end 
          if(!_maxi_write_data_busy && !_maxi_write_req_fifo_empty && (_maxi_write_op_sel_fifo == 2)) begin
            _maxi_write_data_fsm <= _maxi_write_data_fsm_1;
          end 
          if(!_maxi_write_data_busy && !_maxi_write_req_fifo_empty && (_maxi_write_op_sel_fifo == 3)) begin
            _maxi_write_data_fsm <= _maxi_write_data_fsm_1;
          end 
        end
        _maxi_write_data_fsm_1: begin
          _maxi_write_data_fsm <= _maxi_write_data_fsm_2;
          _maxi_write_data_fsm <= _maxi_write_data_fsm_2;
          _maxi_write_data_fsm <= _maxi_write_data_fsm_2;
        end
        _maxi_write_data_fsm_2: begin
          if((_maxi_write_op_sel_buf == 1) && read_burst_packed_rvalid_1308 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)) && read_burst_packed_rlast_1309) begin
            _maxi_write_data_fsm <= _maxi_write_data_fsm_init;
          end 
          if((_maxi_write_op_sel_buf == 2) && read_burst_packed_rvalid_1456 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)) && read_burst_packed_rlast_1457) begin
            _maxi_write_data_fsm <= _maxi_write_data_fsm_init;
          end 
          if((_maxi_write_op_sel_buf == 3) && read_burst_packed_rvalid_1608 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)) && read_burst_packed_rlast_1609) begin
            _maxi_write_data_fsm <= _maxi_write_data_fsm_init;
          end 
        end
      endcase
    end
  end

  localparam read_burst_packed_fsm_24_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      read_burst_packed_fsm_24 <= read_burst_packed_fsm_24_init;
      read_burst_packed_addr_1305 <= 0;
      read_burst_packed_stride_1306 <= 0;
      read_burst_packed_length_1307 <= 0;
      read_burst_packed_rvalid_1308 <= 0;
      read_burst_packed_rlast_1309 <= 0;
    end else begin
      case(read_burst_packed_fsm_24)
        read_burst_packed_fsm_24_init: begin
          read_burst_packed_addr_1305 <= _maxi_write_local_addr_buf;
          read_burst_packed_stride_1306 <= _maxi_write_local_stride_buf;
          read_burst_packed_length_1307 <= _maxi_write_size_buf;
          read_burst_packed_rvalid_1308 <= 0;
          read_burst_packed_rlast_1309 <= 0;
          if((_maxi_write_data_fsm == 1) && (_maxi_write_op_sel_buf == 1) && (_maxi_write_size_buf > 0)) begin
            read_burst_packed_fsm_24 <= read_burst_packed_fsm_24_1;
          end 
        end
        read_burst_packed_fsm_24_1: begin
          if((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0) && (read_burst_packed_length_1307 > 0)) begin
            read_burst_packed_addr_1305 <= read_burst_packed_addr_1305 + read_burst_packed_stride_1306;
            read_burst_packed_length_1307 <= read_burst_packed_length_1307 - 1;
            read_burst_packed_rvalid_1308 <= 1;
          end 
          if((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0) && (read_burst_packed_length_1307 <= 1)) begin
            read_burst_packed_rlast_1309 <= 1;
          end 
          if(read_burst_packed_rlast_1309 && read_burst_packed_rvalid_1308 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) begin
            read_burst_packed_rvalid_1308 <= 0;
            read_burst_packed_rlast_1309 <= 0;
          end 
          if(0) begin
            read_burst_packed_rvalid_1308 <= 0;
            read_burst_packed_rlast_1309 <= 0;
          end 
          if(read_burst_packed_rlast_1309 && read_burst_packed_rvalid_1308 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) begin
            read_burst_packed_fsm_24 <= read_burst_packed_fsm_24_init;
          end 
          if(0) begin
            read_burst_packed_fsm_24 <= read_burst_packed_fsm_24_init;
          end 
        end
      endcase
    end
  end

  localparam control_max_pool_serial_26_1 = 1;
  localparam control_max_pool_serial_26_2 = 2;
  localparam control_max_pool_serial_26_3 = 3;
  localparam control_max_pool_serial_26_4 = 4;
  localparam control_max_pool_serial_26_5 = 5;
  localparam control_max_pool_serial_26_6 = 6;
  localparam control_max_pool_serial_26_7 = 7;
  localparam control_max_pool_serial_26_8 = 8;
  localparam control_max_pool_serial_26_9 = 9;
  localparam control_max_pool_serial_26_10 = 10;
  localparam control_max_pool_serial_26_11 = 11;
  localparam control_max_pool_serial_26_12 = 12;
  localparam control_max_pool_serial_26_13 = 13;
  localparam control_max_pool_serial_26_14 = 14;
  localparam control_max_pool_serial_26_15 = 15;
  localparam control_max_pool_serial_26_16 = 16;
  localparam control_max_pool_serial_26_17 = 17;
  localparam control_max_pool_serial_26_18 = 18;
  localparam control_max_pool_serial_26_19 = 19;

  always @(posedge CLK) begin
    if(RST) begin
      control_max_pool_serial_26 <= control_max_pool_serial_26_init;
      _control_max_pool_serial_26_called <= 0;
      max_pool_serial_26_act_base_offset_row <= 0;
      max_pool_serial_26_act_base_offset_bat <= 0;
      max_pool_serial_26_act_page <= 0;
      max_pool_serial_26_act_page_comp_offset <= 0;
      max_pool_serial_26_act_page_dma_offset <= 0;
      max_pool_serial_26_out_base_offset_row <= 0;
      max_pool_serial_26_out_base_offset_bat <= 0;
      max_pool_serial_26_out_page <= 0;
      max_pool_serial_26_out_page_comp_offset <= 0;
      max_pool_serial_26_out_page_dma_offset <= 0;
      max_pool_serial_26_row_count <= 0;
      max_pool_serial_26_bat_count <= 0;
      max_pool_serial_26_prev_row_count <= 0;
      max_pool_serial_26_prev_bat_count <= 0;
      max_pool_serial_26_skip_read_act <= 0;
      max_pool_serial_26_skip_comp <= 0;
      max_pool_serial_26_skip_write_out <= 0;
      max_pool_serial_26_out_count <= 0;
    end else begin
      case(control_max_pool_serial_26)
        control_max_pool_serial_26_init: begin
          if(main_fsm == 18) begin
            _control_max_pool_serial_26_called <= 1;
          end 
          if(main_fsm == 35) begin
            _control_max_pool_serial_26_called <= 1;
          end 
          if(main_fsm == 62) begin
            _control_max_pool_serial_26_called <= 1;
          end 
          if(main_fsm == 89) begin
            _control_max_pool_serial_26_called <= 1;
          end 
          if(main_fsm == 116) begin
            _control_max_pool_serial_26_called <= 1;
          end 
          if(main_fsm == 18) begin
            control_max_pool_serial_26 <= control_max_pool_serial_26_1;
          end 
          if(main_fsm == 35) begin
            control_max_pool_serial_26 <= control_max_pool_serial_26_1;
          end 
          if(main_fsm == 62) begin
            control_max_pool_serial_26 <= control_max_pool_serial_26_1;
          end 
          if(main_fsm == 89) begin
            control_max_pool_serial_26 <= control_max_pool_serial_26_1;
          end 
          if(main_fsm == 116) begin
            control_max_pool_serial_26 <= control_max_pool_serial_26_1;
          end 
        end
        control_max_pool_serial_26_1: begin
          control_max_pool_serial_26 <= control_max_pool_serial_26_2;
        end
        control_max_pool_serial_26_2: begin
          max_pool_serial_26_act_base_offset_row <= 0;
          max_pool_serial_26_act_base_offset_bat <= 0;
          max_pool_serial_26_act_page <= 0;
          max_pool_serial_26_act_page_comp_offset <= 0;
          max_pool_serial_26_act_page_dma_offset <= 0;
          max_pool_serial_26_out_base_offset_row <= 0;
          max_pool_serial_26_out_base_offset_bat <= 0;
          max_pool_serial_26_out_page <= 0;
          max_pool_serial_26_out_page_comp_offset <= 0;
          max_pool_serial_26_out_page_dma_offset <= 0;
          max_pool_serial_26_row_count <= 0;
          max_pool_serial_26_bat_count <= 0;
          max_pool_serial_26_prev_row_count <= 0;
          max_pool_serial_26_prev_bat_count <= 0;
          max_pool_serial_26_skip_read_act <= 0;
          max_pool_serial_26_skip_comp <= 0;
          max_pool_serial_26_skip_write_out <= 1;
          max_pool_serial_26_out_count <= 0;
          control_max_pool_serial_26 <= control_max_pool_serial_26_3;
        end
        control_max_pool_serial_26_3: begin
          control_max_pool_serial_26 <= control_max_pool_serial_26_4;
          if(max_pool_serial_26_skip_read_act) begin
            control_max_pool_serial_26 <= control_max_pool_serial_26_11;
          end 
        end
        control_max_pool_serial_26_4: begin
          control_max_pool_serial_26 <= control_max_pool_serial_26_5;
          if(max_pool_serial_26_dma_pad_mask_0) begin
            control_max_pool_serial_26 <= control_max_pool_serial_26_7;
          end 
        end
        control_max_pool_serial_26_5: begin
          if(_maxi_read_req_idle) begin
            control_max_pool_serial_26 <= control_max_pool_serial_26_6;
          end 
        end
        control_max_pool_serial_26_6: begin
          if(_maxi_read_idle) begin
            control_max_pool_serial_26 <= control_max_pool_serial_26_7;
          end 
        end
        control_max_pool_serial_26_7: begin
          control_max_pool_serial_26 <= control_max_pool_serial_26_8;
          if(max_pool_serial_26_dma_pad_mask_1) begin
            control_max_pool_serial_26 <= control_max_pool_serial_26_10;
          end 
        end
        control_max_pool_serial_26_8: begin
          if(_maxi_read_req_idle) begin
            control_max_pool_serial_26 <= control_max_pool_serial_26_9;
          end 
        end
        control_max_pool_serial_26_9: begin
          if(_maxi_read_idle) begin
            control_max_pool_serial_26 <= control_max_pool_serial_26_10;
          end 
        end
        control_max_pool_serial_26_10: begin
          control_max_pool_serial_26 <= control_max_pool_serial_26_11;
        end
        control_max_pool_serial_26_11: begin
          if(_maxi_write_idle) begin
            control_max_pool_serial_26 <= control_max_pool_serial_26_12;
          end 
        end
        control_max_pool_serial_26_12: begin
          if(max_pool_serial_26_comp_fsm == 0) begin
            control_max_pool_serial_26 <= control_max_pool_serial_26_13;
          end 
        end
        control_max_pool_serial_26_13: begin
          control_max_pool_serial_26 <= control_max_pool_serial_26_14;
          if(max_pool_serial_26_skip_write_out) begin
            control_max_pool_serial_26 <= control_max_pool_serial_26_17;
          end 
        end
        control_max_pool_serial_26_14: begin
          if(max_pool_serial_26_comp_count >= max_pool_serial_26_out_count + cparam_max_pool_serial_26_out_write_size) begin
            control_max_pool_serial_26 <= control_max_pool_serial_26_15;
          end 
        end
        control_max_pool_serial_26_15: begin
          if(_maxi_write_req_idle) begin
            control_max_pool_serial_26 <= control_max_pool_serial_26_16;
          end 
        end
        control_max_pool_serial_26_16: begin
          max_pool_serial_26_out_count <= max_pool_serial_26_out_count + cparam_max_pool_serial_26_out_write_size;
          control_max_pool_serial_26 <= control_max_pool_serial_26_17;
        end
        control_max_pool_serial_26_17: begin
          max_pool_serial_26_act_base_offset_row <= max_pool_serial_26_act_base_offset_row + cparam_max_pool_serial_26_act_row_step;
          if(max_pool_serial_26_row_count >= cparam_max_pool_serial_26_max_row_count) begin
            max_pool_serial_26_act_base_offset_row <= 0;
            max_pool_serial_26_act_base_offset_bat <= max_pool_serial_26_act_base_offset_bat + cparam_max_pool_serial_26_act_bat_step;
          end 
          if((max_pool_serial_26_row_count >= cparam_max_pool_serial_26_max_row_count) && (max_pool_serial_26_bat_count >= cparam_max_pool_serial_26_max_bat_count)) begin
            max_pool_serial_26_act_base_offset_bat <= 0;
          end 
          max_pool_serial_26_row_count <= max_pool_serial_26_row_count + cparam_max_pool_serial_26_stride_row;
          if(max_pool_serial_26_row_count >= cparam_max_pool_serial_26_max_row_count) begin
            max_pool_serial_26_row_count <= 0;
            max_pool_serial_26_bat_count <= max_pool_serial_26_bat_count + 1;
          end 
          if((max_pool_serial_26_row_count >= cparam_max_pool_serial_26_max_row_count) && (max_pool_serial_26_bat_count >= cparam_max_pool_serial_26_max_bat_count)) begin
            max_pool_serial_26_bat_count <= 0;
          end 
          if(!max_pool_serial_26_act_page) begin
            max_pool_serial_26_act_page_comp_offset <= 131072;
            max_pool_serial_26_act_page_dma_offset <= 131072;
            max_pool_serial_26_act_page <= 1;
          end 
          if(max_pool_serial_26_act_page) begin
            max_pool_serial_26_act_page_comp_offset <= 0;
            max_pool_serial_26_act_page_dma_offset <= 0;
            max_pool_serial_26_act_page <= 0;
          end 
          if(!max_pool_serial_26_skip_write_out) begin
            max_pool_serial_26_out_base_offset_row <= max_pool_serial_26_out_base_offset_row + cparam_max_pool_serial_26_out_row_step;
          end 
          if(!max_pool_serial_26_skip_write_out && (max_pool_serial_26_prev_row_count >= cparam_max_pool_serial_26_max_row_count)) begin
            max_pool_serial_26_out_base_offset_row <= 0;
            max_pool_serial_26_out_base_offset_bat <= max_pool_serial_26_out_base_offset_bat + cparam_max_pool_serial_26_out_bat_step;
          end 
          if(!max_pool_serial_26_skip_write_out && (max_pool_serial_26_prev_row_count >= cparam_max_pool_serial_26_max_row_count) && (max_pool_serial_26_prev_bat_count >= cparam_max_pool_serial_26_max_bat_count)) begin
            max_pool_serial_26_out_base_offset_bat <= 0;
          end 
          if(!max_pool_serial_26_out_page) begin
            max_pool_serial_26_out_page_comp_offset <= 8192;
            max_pool_serial_26_out_page_dma_offset <= 0;
            max_pool_serial_26_out_page <= 1;
          end 
          if(max_pool_serial_26_out_page) begin
            max_pool_serial_26_out_page_comp_offset <= 0;
            max_pool_serial_26_out_page_dma_offset <= 8192;
            max_pool_serial_26_out_page <= 0;
          end 
          max_pool_serial_26_prev_row_count <= max_pool_serial_26_row_count;
          max_pool_serial_26_prev_bat_count <= max_pool_serial_26_bat_count;
          if((max_pool_serial_26_row_count >= cparam_max_pool_serial_26_max_row_count) && (max_pool_serial_26_bat_count >= cparam_max_pool_serial_26_max_bat_count)) begin
            max_pool_serial_26_skip_read_act <= 1;
          end 
          if((max_pool_serial_26_row_count >= cparam_max_pool_serial_26_max_row_count) && (max_pool_serial_26_bat_count >= cparam_max_pool_serial_26_max_bat_count)) begin
            max_pool_serial_26_skip_comp <= 1;
          end 
          if(max_pool_serial_26_skip_write_out && (max_pool_serial_26_prev_row_count == 0) && (max_pool_serial_26_prev_bat_count == 0)) begin
            max_pool_serial_26_skip_write_out <= 0;
          end 
          control_max_pool_serial_26 <= control_max_pool_serial_26_3;
          if(!max_pool_serial_26_skip_write_out && (max_pool_serial_26_prev_row_count >= cparam_max_pool_serial_26_max_row_count) && (max_pool_serial_26_prev_bat_count >= cparam_max_pool_serial_26_max_bat_count)) begin
            control_max_pool_serial_26 <= control_max_pool_serial_26_18;
          end 
        end
        control_max_pool_serial_26_18: begin
          if(_maxi_write_idle && !_maxi_has_outstanding_write) begin
            control_max_pool_serial_26 <= control_max_pool_serial_26_19;
          end 
        end
        control_max_pool_serial_26_19: begin
          if(main_fsm == 21) begin
            _control_max_pool_serial_26_called <= 0;
          end 
          if(main_fsm == 38) begin
            _control_max_pool_serial_26_called <= 0;
          end 
          if(main_fsm == 65) begin
            _control_max_pool_serial_26_called <= 0;
          end 
          if(main_fsm == 92) begin
            _control_max_pool_serial_26_called <= 0;
          end 
          if(main_fsm == 119) begin
            _control_max_pool_serial_26_called <= 0;
          end 
          if(main_fsm == 21) begin
            control_max_pool_serial_26 <= control_max_pool_serial_26_init;
          end 
          if(main_fsm == 38) begin
            control_max_pool_serial_26 <= control_max_pool_serial_26_init;
          end 
          if(main_fsm == 65) begin
            control_max_pool_serial_26 <= control_max_pool_serial_26_init;
          end 
          if(main_fsm == 92) begin
            control_max_pool_serial_26 <= control_max_pool_serial_26_init;
          end 
          if(main_fsm == 119) begin
            control_max_pool_serial_26 <= control_max_pool_serial_26_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_25_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_25 <= write_burst_packed_fsm_25_init;
      write_burst_packed_addr_1332 <= 0;
      write_burst_packed_stride_1333 <= 0;
      write_burst_packed_length_1334 <= 0;
      write_burst_packed_done_1335 <= 0;
    end else begin
      case(write_burst_packed_fsm_25)
        write_burst_packed_fsm_25_init: begin
          write_burst_packed_addr_1332 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_1333 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_1334 <= _maxi_read_local_size_buf;
          write_burst_packed_done_1335 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 7) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_25 <= write_burst_packed_fsm_25_1;
          end 
        end
        write_burst_packed_fsm_25_1: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_packed_addr_1332 <= write_burst_packed_addr_1332 + write_burst_packed_stride_1333;
            write_burst_packed_length_1334 <= write_burst_packed_length_1334 - 1;
            write_burst_packed_done_1335 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_packed_length_1334 <= 1)) begin
            write_burst_packed_done_1335 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_packed_done_1335 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_packed_length_1334 <= 1)) begin
            write_burst_packed_fsm_25 <= write_burst_packed_fsm_25_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_packed_fsm_25 <= write_burst_packed_fsm_25_init;
          end 
          if(0) begin
            write_burst_packed_fsm_25 <= write_burst_packed_fsm_25_init;
          end 
        end
      endcase
    end
  end

  localparam max_pool_serial_26_comp_fsm_1 = 1;
  localparam max_pool_serial_26_comp_fsm_2 = 2;
  localparam max_pool_serial_26_comp_fsm_3 = 3;
  localparam max_pool_serial_26_comp_fsm_4 = 4;
  localparam max_pool_serial_26_comp_fsm_5 = 5;
  localparam max_pool_serial_26_comp_fsm_6 = 6;
  localparam max_pool_serial_26_comp_fsm_7 = 7;

  always @(posedge CLK) begin
    if(RST) begin
      max_pool_serial_26_comp_fsm <= max_pool_serial_26_comp_fsm_init;
      max_pool_serial_26_stream_act_local <= 0;
      max_pool_serial_26_stream_out_local <= 0;
      max_pool_serial_26_col_count <= 0;
      max_pool_serial_26_act_page_comp_offset_buf <= 0;
      max_pool_serial_26_out_page_comp_offset_buf <= 0;
      max_pool_serial_26_row_count_buf <= 0;
      max_pool_serial_26_stream_pad_masks <= 0;
      max_pool_serial_26_comp_count <= 0;
    end else begin
      if(control_max_pool_serial_26 == 2) begin
        max_pool_serial_26_comp_count <= 0;
      end 
      if(_stream_max_pool_serial_26_sink_stop) begin
        max_pool_serial_26_comp_count <= max_pool_serial_26_comp_count + cparam_max_pool_serial_26_inc_out_laddr;
      end 
      case(max_pool_serial_26_comp_fsm)
        max_pool_serial_26_comp_fsm_init: begin
          if((control_max_pool_serial_26 == 12) && !max_pool_serial_26_skip_comp) begin
            max_pool_serial_26_comp_fsm <= max_pool_serial_26_comp_fsm_1;
          end 
        end
        max_pool_serial_26_comp_fsm_1: begin
          max_pool_serial_26_stream_act_local <= cparam_max_pool_serial_26_local_pad_offset;
          max_pool_serial_26_stream_out_local <= 0;
          max_pool_serial_26_col_count <= 0;
          max_pool_serial_26_act_page_comp_offset_buf <= max_pool_serial_26_act_page_comp_offset;
          max_pool_serial_26_out_page_comp_offset_buf <= max_pool_serial_26_out_page_comp_offset;
          max_pool_serial_26_row_count_buf <= max_pool_serial_26_row_count;
          max_pool_serial_26_comp_fsm <= max_pool_serial_26_comp_fsm_2;
        end
        max_pool_serial_26_comp_fsm_2: begin
          max_pool_serial_26_stream_pad_masks <= { max_pool_serial_26_stream_pad_mask_1_1, max_pool_serial_26_stream_pad_mask_1_0, max_pool_serial_26_stream_pad_mask_0_1, max_pool_serial_26_stream_pad_mask_0_0 };
          max_pool_serial_26_comp_fsm <= max_pool_serial_26_comp_fsm_3;
        end
        max_pool_serial_26_comp_fsm_3: begin
          if(!_stream_max_pool_serial_26_source_busy) begin
            max_pool_serial_26_comp_fsm <= max_pool_serial_26_comp_fsm_4;
          end 
        end
        max_pool_serial_26_comp_fsm_4: begin
          max_pool_serial_26_comp_fsm <= max_pool_serial_26_comp_fsm_5;
          max_pool_serial_26_comp_fsm <= max_pool_serial_26_comp_fsm_5;
          max_pool_serial_26_comp_fsm <= max_pool_serial_26_comp_fsm_5;
          if(_stream_max_pool_serial_26_stream_oready) begin
            max_pool_serial_26_comp_fsm <= max_pool_serial_26_comp_fsm_5;
          end 
        end
        max_pool_serial_26_comp_fsm_5: begin
          max_pool_serial_26_comp_fsm <= max_pool_serial_26_comp_fsm_6;
        end
        max_pool_serial_26_comp_fsm_6: begin
          if(_stream_max_pool_serial_26_busy) begin
            max_pool_serial_26_comp_fsm <= max_pool_serial_26_comp_fsm_7;
          end 
        end
        max_pool_serial_26_comp_fsm_7: begin
          max_pool_serial_26_stream_act_local <= max_pool_serial_26_stream_act_local + cparam_max_pool_serial_26_inc_act_laddr;
          if(max_pool_serial_26_col_count >= cparam_max_pool_serial_26_max_col_count) begin
            max_pool_serial_26_stream_act_local <= cparam_max_pool_serial_26_local_pad_offset;
          end 
          max_pool_serial_26_stream_out_local <= max_pool_serial_26_stream_out_local + cparam_max_pool_serial_26_inc_out_laddr;
          if(max_pool_serial_26_col_count >= cparam_max_pool_serial_26_max_col_count) begin
            max_pool_serial_26_stream_out_local <= 0;
          end 
          max_pool_serial_26_col_count <= max_pool_serial_26_col_count + cparam_max_pool_serial_26_stride_col;
          if(max_pool_serial_26_col_count >= cparam_max_pool_serial_26_max_col_count) begin
            max_pool_serial_26_col_count <= 0;
          end 
          max_pool_serial_26_comp_fsm <= max_pool_serial_26_comp_fsm_2;
          if(max_pool_serial_26_col_count >= cparam_max_pool_serial_26_max_col_count) begin
            max_pool_serial_26_comp_fsm <= max_pool_serial_26_comp_fsm_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_1353 <= 0;
      _tmp_1704 <= 0;
    end else begin
      if(_stream_max_pool_serial_26_stream_oready && _stream_max_pool_serial_26_source_1_source_ram_renable && (_stream_max_pool_serial_26_source_1_source_sel == 1)) begin
        _tmp_1353 <= read_rtl_bank_1352;
      end 
      if(_stream_matmul_55_stream_oready && _stream_matmul_55_source_21_source_ram_renable && (_stream_matmul_55_source_21_source_sel == 4)) begin
        _tmp_1704 <= read_rtl_bank_1703;
      end 
    end
  end

  localparam _stream_max_pool_serial_26_source_1_source_pat_fsm_0_1 = 1;
  localparam _stream_max_pool_serial_26_source_1_source_pat_fsm_0_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_max_pool_serial_26_source_1_source_pat_fsm_0 <= _stream_max_pool_serial_26_source_1_source_pat_fsm_0_init;
    end else begin
      case(_stream_max_pool_serial_26_source_1_source_pat_fsm_0)
        _stream_max_pool_serial_26_source_1_source_pat_fsm_0_init: begin
          if(_stream_max_pool_serial_26_source_start && _stream_max_pool_serial_26_source_1_source_mode & 5'b10 && _stream_max_pool_serial_26_stream_oready) begin
            _stream_max_pool_serial_26_source_1_source_pat_fsm_0 <= _stream_max_pool_serial_26_source_1_source_pat_fsm_0_1;
          end 
        end
        _stream_max_pool_serial_26_source_1_source_pat_fsm_0_1: begin
          if(_stream_max_pool_serial_26_source_stop && _stream_max_pool_serial_26_stream_oready) begin
            _stream_max_pool_serial_26_source_1_source_pat_fsm_0 <= _stream_max_pool_serial_26_source_1_source_pat_fsm_0_init;
          end 
          if((_source_stream_max_pool_serial_26_source_1_pat_count_0 == 0) && (_source_stream_max_pool_serial_26_source_1_pat_count_1 == 0) && (_source_stream_max_pool_serial_26_source_1_pat_count_2 == 0) && (_source_stream_max_pool_serial_26_source_1_pat_count_3 == 0) && _stream_max_pool_serial_26_stream_oready) begin
            _stream_max_pool_serial_26_source_1_source_pat_fsm_0 <= _stream_max_pool_serial_26_source_1_source_pat_fsm_0_2;
          end 
        end
        _stream_max_pool_serial_26_source_1_source_pat_fsm_0_2: begin
          if(_stream_max_pool_serial_26_stream_oready) begin
            _stream_max_pool_serial_26_source_1_source_pat_fsm_0 <= _stream_max_pool_serial_26_source_1_source_pat_fsm_0_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_max_pool_serial_26_sink_5_sink_fsm_1_1 = 1;
  localparam _stream_max_pool_serial_26_sink_5_sink_fsm_1_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_max_pool_serial_26_sink_5_sink_fsm_1 <= _stream_max_pool_serial_26_sink_5_sink_fsm_1_init;
    end else begin
      case(_stream_max_pool_serial_26_sink_5_sink_fsm_1)
        _stream_max_pool_serial_26_sink_5_sink_fsm_1_init: begin
          if(_stream_max_pool_serial_26_sink_start && _stream_max_pool_serial_26_sink_5_sink_mode & 5'b1 && _stream_max_pool_serial_26_stream_oready) begin
            _stream_max_pool_serial_26_sink_5_sink_fsm_1 <= _stream_max_pool_serial_26_sink_5_sink_fsm_1_1;
          end 
        end
        _stream_max_pool_serial_26_sink_5_sink_fsm_1_1: begin
          if(_stream_max_pool_serial_26_stream_oready) begin
            _stream_max_pool_serial_26_sink_5_sink_fsm_1 <= _stream_max_pool_serial_26_sink_5_sink_fsm_1_2;
          end 
        end
        _stream_max_pool_serial_26_sink_5_sink_fsm_1_2: begin
          if(stream_max_pool_serial_26_sink_6_data && (_stream_max_pool_serial_26_sink_5_sink_count == 1) && _stream_max_pool_serial_26_stream_oready) begin
            _stream_max_pool_serial_26_sink_5_sink_fsm_1 <= _stream_max_pool_serial_26_sink_5_sink_fsm_1_init;
          end 
          if(_stream_max_pool_serial_26_sink_stop && _stream_max_pool_serial_26_stream_oready) begin
            _stream_max_pool_serial_26_sink_5_sink_fsm_1 <= _stream_max_pool_serial_26_sink_5_sink_fsm_1_init;
          end 
        end
      endcase
    end
  end

  localparam read_burst_packed_fsm_26_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      read_burst_packed_fsm_26 <= read_burst_packed_fsm_26_init;
      read_burst_packed_addr_1453 <= 0;
      read_burst_packed_stride_1454 <= 0;
      read_burst_packed_length_1455 <= 0;
      read_burst_packed_rvalid_1456 <= 0;
      read_burst_packed_rlast_1457 <= 0;
    end else begin
      case(read_burst_packed_fsm_26)
        read_burst_packed_fsm_26_init: begin
          read_burst_packed_addr_1453 <= _maxi_write_local_addr_buf;
          read_burst_packed_stride_1454 <= _maxi_write_local_stride_buf;
          read_burst_packed_length_1455 <= _maxi_write_size_buf;
          read_burst_packed_rvalid_1456 <= 0;
          read_burst_packed_rlast_1457 <= 0;
          if((_maxi_write_data_fsm == 1) && (_maxi_write_op_sel_buf == 2) && (_maxi_write_size_buf > 0)) begin
            read_burst_packed_fsm_26 <= read_burst_packed_fsm_26_1;
          end 
        end
        read_burst_packed_fsm_26_1: begin
          if((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0) && (read_burst_packed_length_1455 > 0)) begin
            read_burst_packed_addr_1453 <= read_burst_packed_addr_1453 + read_burst_packed_stride_1454;
            read_burst_packed_length_1455 <= read_burst_packed_length_1455 - 1;
            read_burst_packed_rvalid_1456 <= 1;
          end 
          if((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0) && (read_burst_packed_length_1455 <= 1)) begin
            read_burst_packed_rlast_1457 <= 1;
          end 
          if(read_burst_packed_rlast_1457 && read_burst_packed_rvalid_1456 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) begin
            read_burst_packed_rvalid_1456 <= 0;
            read_burst_packed_rlast_1457 <= 0;
          end 
          if(0) begin
            read_burst_packed_rvalid_1456 <= 0;
            read_burst_packed_rlast_1457 <= 0;
          end 
          if(read_burst_packed_rlast_1457 && read_burst_packed_rvalid_1456 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) begin
            read_burst_packed_fsm_26 <= read_burst_packed_fsm_26_init;
          end 
          if(0) begin
            read_burst_packed_fsm_26 <= read_burst_packed_fsm_26_init;
          end 
        end
      endcase
    end
  end

  localparam control_avg_pool_serial_52_1 = 1;
  localparam control_avg_pool_serial_52_2 = 2;
  localparam control_avg_pool_serial_52_3 = 3;
  localparam control_avg_pool_serial_52_4 = 4;
  localparam control_avg_pool_serial_52_5 = 5;
  localparam control_avg_pool_serial_52_6 = 6;
  localparam control_avg_pool_serial_52_7 = 7;
  localparam control_avg_pool_serial_52_8 = 8;
  localparam control_avg_pool_serial_52_9 = 9;
  localparam control_avg_pool_serial_52_10 = 10;
  localparam control_avg_pool_serial_52_11 = 11;
  localparam control_avg_pool_serial_52_12 = 12;
  localparam control_avg_pool_serial_52_13 = 13;
  localparam control_avg_pool_serial_52_14 = 14;
  localparam control_avg_pool_serial_52_15 = 15;
  localparam control_avg_pool_serial_52_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      control_avg_pool_serial_52 <= control_avg_pool_serial_52_init;
      _control_avg_pool_serial_52_called <= 0;
      avg_pool_serial_52_act_base_offset_row <= 0;
      avg_pool_serial_52_act_base_offset_bat <= 0;
      avg_pool_serial_52_act_page <= 0;
      avg_pool_serial_52_act_page_comp_offset <= 0;
      avg_pool_serial_52_act_page_dma_offset <= 0;
      avg_pool_serial_52_out_base_offset_row <= 0;
      avg_pool_serial_52_out_base_offset_bat <= 0;
      avg_pool_serial_52_out_page <= 0;
      avg_pool_serial_52_out_page_comp_offset <= 0;
      avg_pool_serial_52_out_page_dma_offset <= 0;
      avg_pool_serial_52_row_count <= 0;
      avg_pool_serial_52_bat_count <= 0;
      avg_pool_serial_52_prev_row_count <= 0;
      avg_pool_serial_52_prev_bat_count <= 0;
      avg_pool_serial_52_skip_read_act <= 0;
      avg_pool_serial_52_skip_comp <= 0;
      avg_pool_serial_52_skip_write_out <= 0;
      avg_pool_serial_52_out_count <= 0;
    end else begin
      case(control_avg_pool_serial_52)
        control_avg_pool_serial_52_init: begin
          if(main_fsm == 122) begin
            _control_avg_pool_serial_52_called <= 1;
          end 
          if(main_fsm == 122) begin
            control_avg_pool_serial_52 <= control_avg_pool_serial_52_1;
          end 
        end
        control_avg_pool_serial_52_1: begin
          control_avg_pool_serial_52 <= control_avg_pool_serial_52_2;
        end
        control_avg_pool_serial_52_2: begin
          avg_pool_serial_52_act_base_offset_row <= 0;
          avg_pool_serial_52_act_base_offset_bat <= 0;
          avg_pool_serial_52_act_page <= 0;
          avg_pool_serial_52_act_page_comp_offset <= 0;
          avg_pool_serial_52_act_page_dma_offset <= 0;
          avg_pool_serial_52_out_base_offset_row <= 0;
          avg_pool_serial_52_out_base_offset_bat <= 0;
          avg_pool_serial_52_out_page <= 0;
          avg_pool_serial_52_out_page_comp_offset <= 0;
          avg_pool_serial_52_out_page_dma_offset <= 0;
          avg_pool_serial_52_row_count <= 0;
          avg_pool_serial_52_bat_count <= 0;
          avg_pool_serial_52_prev_row_count <= 0;
          avg_pool_serial_52_prev_bat_count <= 0;
          avg_pool_serial_52_skip_read_act <= 0;
          avg_pool_serial_52_skip_comp <= 0;
          avg_pool_serial_52_skip_write_out <= 1;
          avg_pool_serial_52_out_count <= 0;
          control_avg_pool_serial_52 <= control_avg_pool_serial_52_3;
        end
        control_avg_pool_serial_52_3: begin
          control_avg_pool_serial_52 <= control_avg_pool_serial_52_4;
          if(avg_pool_serial_52_skip_read_act) begin
            control_avg_pool_serial_52 <= control_avg_pool_serial_52_8;
          end 
        end
        control_avg_pool_serial_52_4: begin
          control_avg_pool_serial_52 <= control_avg_pool_serial_52_5;
          if(avg_pool_serial_52_dma_pad_mask_0) begin
            control_avg_pool_serial_52 <= control_avg_pool_serial_52_7;
          end 
        end
        control_avg_pool_serial_52_5: begin
          if(_maxi_read_req_idle) begin
            control_avg_pool_serial_52 <= control_avg_pool_serial_52_6;
          end 
        end
        control_avg_pool_serial_52_6: begin
          if(_maxi_read_idle) begin
            control_avg_pool_serial_52 <= control_avg_pool_serial_52_7;
          end 
        end
        control_avg_pool_serial_52_7: begin
          control_avg_pool_serial_52 <= control_avg_pool_serial_52_8;
        end
        control_avg_pool_serial_52_8: begin
          if(_maxi_write_idle) begin
            control_avg_pool_serial_52 <= control_avg_pool_serial_52_9;
          end 
        end
        control_avg_pool_serial_52_9: begin
          if(avg_pool_serial_52_comp_fsm == 0) begin
            control_avg_pool_serial_52 <= control_avg_pool_serial_52_10;
          end 
        end
        control_avg_pool_serial_52_10: begin
          control_avg_pool_serial_52 <= control_avg_pool_serial_52_11;
          if(avg_pool_serial_52_skip_write_out) begin
            control_avg_pool_serial_52 <= control_avg_pool_serial_52_14;
          end 
        end
        control_avg_pool_serial_52_11: begin
          if(avg_pool_serial_52_comp_count >= avg_pool_serial_52_out_count + cparam_avg_pool_serial_52_out_write_size) begin
            control_avg_pool_serial_52 <= control_avg_pool_serial_52_12;
          end 
        end
        control_avg_pool_serial_52_12: begin
          if(_maxi_write_req_idle) begin
            control_avg_pool_serial_52 <= control_avg_pool_serial_52_13;
          end 
        end
        control_avg_pool_serial_52_13: begin
          avg_pool_serial_52_out_count <= avg_pool_serial_52_out_count + cparam_avg_pool_serial_52_out_write_size;
          control_avg_pool_serial_52 <= control_avg_pool_serial_52_14;
        end
        control_avg_pool_serial_52_14: begin
          avg_pool_serial_52_act_base_offset_row <= avg_pool_serial_52_act_base_offset_row + cparam_avg_pool_serial_52_act_row_step;
          if(avg_pool_serial_52_row_count >= cparam_avg_pool_serial_52_max_row_count) begin
            avg_pool_serial_52_act_base_offset_row <= 0;
            avg_pool_serial_52_act_base_offset_bat <= avg_pool_serial_52_act_base_offset_bat + cparam_avg_pool_serial_52_act_bat_step;
          end 
          if((avg_pool_serial_52_row_count >= cparam_avg_pool_serial_52_max_row_count) && (avg_pool_serial_52_bat_count >= cparam_avg_pool_serial_52_max_bat_count)) begin
            avg_pool_serial_52_act_base_offset_bat <= 0;
          end 
          avg_pool_serial_52_row_count <= avg_pool_serial_52_row_count + cparam_avg_pool_serial_52_stride_row;
          if(avg_pool_serial_52_row_count >= cparam_avg_pool_serial_52_max_row_count) begin
            avg_pool_serial_52_row_count <= 0;
            avg_pool_serial_52_bat_count <= avg_pool_serial_52_bat_count + 1;
          end 
          if((avg_pool_serial_52_row_count >= cparam_avg_pool_serial_52_max_row_count) && (avg_pool_serial_52_bat_count >= cparam_avg_pool_serial_52_max_bat_count)) begin
            avg_pool_serial_52_bat_count <= 0;
          end 
          if(!avg_pool_serial_52_act_page) begin
            avg_pool_serial_52_act_page_comp_offset <= 8192;
            avg_pool_serial_52_act_page_dma_offset <= 8192;
            avg_pool_serial_52_act_page <= 1;
          end 
          if(avg_pool_serial_52_act_page) begin
            avg_pool_serial_52_act_page_comp_offset <= 0;
            avg_pool_serial_52_act_page_dma_offset <= 0;
            avg_pool_serial_52_act_page <= 0;
          end 
          if(!avg_pool_serial_52_skip_write_out) begin
            avg_pool_serial_52_out_base_offset_row <= avg_pool_serial_52_out_base_offset_row + cparam_avg_pool_serial_52_out_row_step;
          end 
          if(!avg_pool_serial_52_skip_write_out && (avg_pool_serial_52_prev_row_count >= cparam_avg_pool_serial_52_max_row_count)) begin
            avg_pool_serial_52_out_base_offset_row <= 0;
            avg_pool_serial_52_out_base_offset_bat <= avg_pool_serial_52_out_base_offset_bat + cparam_avg_pool_serial_52_out_bat_step;
          end 
          if(!avg_pool_serial_52_skip_write_out && (avg_pool_serial_52_prev_row_count >= cparam_avg_pool_serial_52_max_row_count) && (avg_pool_serial_52_prev_bat_count >= cparam_avg_pool_serial_52_max_bat_count)) begin
            avg_pool_serial_52_out_base_offset_bat <= 0;
          end 
          if(!avg_pool_serial_52_out_page) begin
            avg_pool_serial_52_out_page_comp_offset <= 8192;
            avg_pool_serial_52_out_page_dma_offset <= 0;
            avg_pool_serial_52_out_page <= 1;
          end 
          if(avg_pool_serial_52_out_page) begin
            avg_pool_serial_52_out_page_comp_offset <= 0;
            avg_pool_serial_52_out_page_dma_offset <= 8192;
            avg_pool_serial_52_out_page <= 0;
          end 
          avg_pool_serial_52_prev_row_count <= avg_pool_serial_52_row_count;
          avg_pool_serial_52_prev_bat_count <= avg_pool_serial_52_bat_count;
          if((avg_pool_serial_52_row_count >= cparam_avg_pool_serial_52_max_row_count) && (avg_pool_serial_52_bat_count >= cparam_avg_pool_serial_52_max_bat_count)) begin
            avg_pool_serial_52_skip_read_act <= 1;
          end 
          if((avg_pool_serial_52_row_count >= cparam_avg_pool_serial_52_max_row_count) && (avg_pool_serial_52_bat_count >= cparam_avg_pool_serial_52_max_bat_count)) begin
            avg_pool_serial_52_skip_comp <= 1;
          end 
          if(avg_pool_serial_52_skip_write_out && (avg_pool_serial_52_prev_row_count == 0) && (avg_pool_serial_52_prev_bat_count == 0)) begin
            avg_pool_serial_52_skip_write_out <= 0;
          end 
          control_avg_pool_serial_52 <= control_avg_pool_serial_52_3;
          if(!avg_pool_serial_52_skip_write_out && (avg_pool_serial_52_prev_row_count >= cparam_avg_pool_serial_52_max_row_count) && (avg_pool_serial_52_prev_bat_count >= cparam_avg_pool_serial_52_max_bat_count)) begin
            control_avg_pool_serial_52 <= control_avg_pool_serial_52_15;
          end 
        end
        control_avg_pool_serial_52_15: begin
          if(_maxi_write_idle && !_maxi_has_outstanding_write) begin
            control_avg_pool_serial_52 <= control_avg_pool_serial_52_16;
          end 
        end
        control_avg_pool_serial_52_16: begin
          if(main_fsm == 125) begin
            _control_avg_pool_serial_52_called <= 0;
          end 
          if(main_fsm == 125) begin
            control_avg_pool_serial_52 <= control_avg_pool_serial_52_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_27_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_27 <= write_burst_packed_fsm_27_init;
      write_burst_packed_addr_1480 <= 0;
      write_burst_packed_stride_1481 <= 0;
      write_burst_packed_length_1482 <= 0;
      write_burst_packed_done_1483 <= 0;
    end else begin
      case(write_burst_packed_fsm_27)
        write_burst_packed_fsm_27_init: begin
          write_burst_packed_addr_1480 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_1481 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_1482 <= _maxi_read_local_size_buf;
          write_burst_packed_done_1483 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 8) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_27 <= write_burst_packed_fsm_27_1;
          end 
        end
        write_burst_packed_fsm_27_1: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_packed_addr_1480 <= write_burst_packed_addr_1480 + write_burst_packed_stride_1481;
            write_burst_packed_length_1482 <= write_burst_packed_length_1482 - 1;
            write_burst_packed_done_1483 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_packed_length_1482 <= 1)) begin
            write_burst_packed_done_1483 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_packed_done_1483 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_packed_length_1482 <= 1)) begin
            write_burst_packed_fsm_27 <= write_burst_packed_fsm_27_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_packed_fsm_27 <= write_burst_packed_fsm_27_init;
          end 
          if(0) begin
            write_burst_packed_fsm_27 <= write_burst_packed_fsm_27_init;
          end 
        end
      endcase
    end
  end

  localparam avg_pool_serial_52_comp_fsm_1 = 1;
  localparam avg_pool_serial_52_comp_fsm_2 = 2;
  localparam avg_pool_serial_52_comp_fsm_3 = 3;
  localparam avg_pool_serial_52_comp_fsm_4 = 4;
  localparam avg_pool_serial_52_comp_fsm_5 = 5;
  localparam avg_pool_serial_52_comp_fsm_6 = 6;
  localparam avg_pool_serial_52_comp_fsm_7 = 7;

  always @(posedge CLK) begin
    if(RST) begin
      avg_pool_serial_52_comp_fsm <= avg_pool_serial_52_comp_fsm_init;
      avg_pool_serial_52_stream_act_local <= 0;
      avg_pool_serial_52_stream_out_local <= 0;
      avg_pool_serial_52_col_count <= 0;
      avg_pool_serial_52_act_page_comp_offset_buf <= 0;
      avg_pool_serial_52_out_page_comp_offset_buf <= 0;
      avg_pool_serial_52_row_count_buf <= 0;
      avg_pool_serial_52_stream_pad_masks <= 0;
      avg_pool_serial_52_comp_count <= 0;
    end else begin
      if(control_avg_pool_serial_52 == 2) begin
        avg_pool_serial_52_comp_count <= 0;
      end 
      if(_stream_avg_pool_serial_52_sink_stop) begin
        avg_pool_serial_52_comp_count <= avg_pool_serial_52_comp_count + cparam_avg_pool_serial_52_inc_out_laddr;
      end 
      case(avg_pool_serial_52_comp_fsm)
        avg_pool_serial_52_comp_fsm_init: begin
          if((control_avg_pool_serial_52 == 9) && !avg_pool_serial_52_skip_comp) begin
            avg_pool_serial_52_comp_fsm <= avg_pool_serial_52_comp_fsm_1;
          end 
        end
        avg_pool_serial_52_comp_fsm_1: begin
          avg_pool_serial_52_stream_act_local <= cparam_avg_pool_serial_52_local_pad_offset;
          avg_pool_serial_52_stream_out_local <= 0;
          avg_pool_serial_52_col_count <= 0;
          avg_pool_serial_52_act_page_comp_offset_buf <= avg_pool_serial_52_act_page_comp_offset;
          avg_pool_serial_52_out_page_comp_offset_buf <= avg_pool_serial_52_out_page_comp_offset;
          avg_pool_serial_52_row_count_buf <= avg_pool_serial_52_row_count;
          avg_pool_serial_52_comp_fsm <= avg_pool_serial_52_comp_fsm_2;
        end
        avg_pool_serial_52_comp_fsm_2: begin
          avg_pool_serial_52_stream_pad_masks <= { avg_pool_serial_52_stream_pad_mask_0_0 };
          avg_pool_serial_52_comp_fsm <= avg_pool_serial_52_comp_fsm_3;
        end
        avg_pool_serial_52_comp_fsm_3: begin
          if(!_stream_avg_pool_serial_52_source_busy) begin
            avg_pool_serial_52_comp_fsm <= avg_pool_serial_52_comp_fsm_4;
          end 
        end
        avg_pool_serial_52_comp_fsm_4: begin
          avg_pool_serial_52_comp_fsm <= avg_pool_serial_52_comp_fsm_5;
          avg_pool_serial_52_comp_fsm <= avg_pool_serial_52_comp_fsm_5;
          avg_pool_serial_52_comp_fsm <= avg_pool_serial_52_comp_fsm_5;
          if(_stream_avg_pool_serial_52_stream_oready) begin
            avg_pool_serial_52_comp_fsm <= avg_pool_serial_52_comp_fsm_5;
          end 
        end
        avg_pool_serial_52_comp_fsm_5: begin
          avg_pool_serial_52_comp_fsm <= avg_pool_serial_52_comp_fsm_6;
        end
        avg_pool_serial_52_comp_fsm_6: begin
          if(_stream_avg_pool_serial_52_busy) begin
            avg_pool_serial_52_comp_fsm <= avg_pool_serial_52_comp_fsm_7;
          end 
        end
        avg_pool_serial_52_comp_fsm_7: begin
          avg_pool_serial_52_stream_act_local <= avg_pool_serial_52_stream_act_local + cparam_avg_pool_serial_52_inc_act_laddr;
          if(avg_pool_serial_52_col_count >= cparam_avg_pool_serial_52_max_col_count) begin
            avg_pool_serial_52_stream_act_local <= cparam_avg_pool_serial_52_local_pad_offset;
          end 
          avg_pool_serial_52_stream_out_local <= avg_pool_serial_52_stream_out_local + cparam_avg_pool_serial_52_inc_out_laddr;
          if(avg_pool_serial_52_col_count >= cparam_avg_pool_serial_52_max_col_count) begin
            avg_pool_serial_52_stream_out_local <= 0;
          end 
          avg_pool_serial_52_col_count <= avg_pool_serial_52_col_count + cparam_avg_pool_serial_52_stride_col;
          if(avg_pool_serial_52_col_count >= cparam_avg_pool_serial_52_max_col_count) begin
            avg_pool_serial_52_col_count <= 0;
          end 
          avg_pool_serial_52_comp_fsm <= avg_pool_serial_52_comp_fsm_2;
          if(avg_pool_serial_52_col_count >= cparam_avg_pool_serial_52_max_col_count) begin
            avg_pool_serial_52_comp_fsm <= avg_pool_serial_52_comp_fsm_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_avg_pool_serial_52_source_1_source_pat_fsm_0_1 = 1;
  localparam _stream_avg_pool_serial_52_source_1_source_pat_fsm_0_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_avg_pool_serial_52_source_1_source_pat_fsm_0 <= _stream_avg_pool_serial_52_source_1_source_pat_fsm_0_init;
    end else begin
      case(_stream_avg_pool_serial_52_source_1_source_pat_fsm_0)
        _stream_avg_pool_serial_52_source_1_source_pat_fsm_0_init: begin
          if(_stream_avg_pool_serial_52_source_start && _stream_avg_pool_serial_52_source_1_source_mode & 5'b10 && _stream_avg_pool_serial_52_stream_oready) begin
            _stream_avg_pool_serial_52_source_1_source_pat_fsm_0 <= _stream_avg_pool_serial_52_source_1_source_pat_fsm_0_1;
          end 
        end
        _stream_avg_pool_serial_52_source_1_source_pat_fsm_0_1: begin
          if(_stream_avg_pool_serial_52_source_stop && _stream_avg_pool_serial_52_stream_oready) begin
            _stream_avg_pool_serial_52_source_1_source_pat_fsm_0 <= _stream_avg_pool_serial_52_source_1_source_pat_fsm_0_init;
          end 
          if((_source_stream_avg_pool_serial_52_source_1_pat_count_0 == 0) && (_source_stream_avg_pool_serial_52_source_1_pat_count_1 == 0) && (_source_stream_avg_pool_serial_52_source_1_pat_count_2 == 0) && (_source_stream_avg_pool_serial_52_source_1_pat_count_3 == 0) && _stream_avg_pool_serial_52_stream_oready) begin
            _stream_avg_pool_serial_52_source_1_source_pat_fsm_0 <= _stream_avg_pool_serial_52_source_1_source_pat_fsm_0_2;
          end 
        end
        _stream_avg_pool_serial_52_source_1_source_pat_fsm_0_2: begin
          if(_stream_avg_pool_serial_52_stream_oready) begin
            _stream_avg_pool_serial_52_source_1_source_pat_fsm_0 <= _stream_avg_pool_serial_52_source_1_source_pat_fsm_0_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_avg_pool_serial_52_sink_5_sink_fsm_1_1 = 1;
  localparam _stream_avg_pool_serial_52_sink_5_sink_fsm_1_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_avg_pool_serial_52_sink_5_sink_fsm_1 <= _stream_avg_pool_serial_52_sink_5_sink_fsm_1_init;
    end else begin
      case(_stream_avg_pool_serial_52_sink_5_sink_fsm_1)
        _stream_avg_pool_serial_52_sink_5_sink_fsm_1_init: begin
          if(_stream_avg_pool_serial_52_sink_start && _stream_avg_pool_serial_52_sink_5_sink_mode & 5'b1 && _stream_avg_pool_serial_52_stream_oready) begin
            _stream_avg_pool_serial_52_sink_5_sink_fsm_1 <= _stream_avg_pool_serial_52_sink_5_sink_fsm_1_1;
          end 
        end
        _stream_avg_pool_serial_52_sink_5_sink_fsm_1_1: begin
          if(_stream_avg_pool_serial_52_stream_oready) begin
            _stream_avg_pool_serial_52_sink_5_sink_fsm_1 <= _stream_avg_pool_serial_52_sink_5_sink_fsm_1_2;
          end 
        end
        _stream_avg_pool_serial_52_sink_5_sink_fsm_1_2: begin
          if(stream_avg_pool_serial_52_sink_6_data && (_stream_avg_pool_serial_52_sink_5_sink_count == 1) && _stream_avg_pool_serial_52_stream_oready) begin
            _stream_avg_pool_serial_52_sink_5_sink_fsm_1 <= _stream_avg_pool_serial_52_sink_5_sink_fsm_1_init;
          end 
          if(_stream_avg_pool_serial_52_sink_stop && _stream_avg_pool_serial_52_stream_oready) begin
            _stream_avg_pool_serial_52_sink_5_sink_fsm_1 <= _stream_avg_pool_serial_52_sink_5_sink_fsm_1_init;
          end 
        end
      endcase
    end
  end

  localparam read_burst_packed_fsm_28_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      read_burst_packed_fsm_28 <= read_burst_packed_fsm_28_init;
      read_burst_packed_addr_1605 <= 0;
      read_burst_packed_stride_1606 <= 0;
      read_burst_packed_length_1607 <= 0;
      read_burst_packed_rvalid_1608 <= 0;
      read_burst_packed_rlast_1609 <= 0;
    end else begin
      case(read_burst_packed_fsm_28)
        read_burst_packed_fsm_28_init: begin
          read_burst_packed_addr_1605 <= _maxi_write_local_addr_buf;
          read_burst_packed_stride_1606 <= _maxi_write_local_stride_buf;
          read_burst_packed_length_1607 <= _maxi_write_size_buf;
          read_burst_packed_rvalid_1608 <= 0;
          read_burst_packed_rlast_1609 <= 0;
          if((_maxi_write_data_fsm == 1) && (_maxi_write_op_sel_buf == 3) && (_maxi_write_size_buf > 0)) begin
            read_burst_packed_fsm_28 <= read_burst_packed_fsm_28_1;
          end 
        end
        read_burst_packed_fsm_28_1: begin
          if((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0) && (read_burst_packed_length_1607 > 0)) begin
            read_burst_packed_addr_1605 <= read_burst_packed_addr_1605 + read_burst_packed_stride_1606;
            read_burst_packed_length_1607 <= read_burst_packed_length_1607 - 1;
            read_burst_packed_rvalid_1608 <= 1;
          end 
          if((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0) && (read_burst_packed_length_1607 <= 1)) begin
            read_burst_packed_rlast_1609 <= 1;
          end 
          if(read_burst_packed_rlast_1609 && read_burst_packed_rvalid_1608 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) begin
            read_burst_packed_rvalid_1608 <= 0;
            read_burst_packed_rlast_1609 <= 0;
          end 
          if(0) begin
            read_burst_packed_rvalid_1608 <= 0;
            read_burst_packed_rlast_1609 <= 0;
          end 
          if(read_burst_packed_rlast_1609 && read_burst_packed_rvalid_1608 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) begin
            read_burst_packed_fsm_28 <= read_burst_packed_fsm_28_init;
          end 
          if(0) begin
            read_burst_packed_fsm_28 <= read_burst_packed_fsm_28_init;
          end 
        end
      endcase
    end
  end

  localparam control_matmul_55_1 = 1;
  localparam control_matmul_55_2 = 2;
  localparam control_matmul_55_3 = 3;
  localparam control_matmul_55_4 = 4;
  localparam control_matmul_55_5 = 5;
  localparam control_matmul_55_6 = 6;
  localparam control_matmul_55_7 = 7;
  localparam control_matmul_55_8 = 8;
  localparam control_matmul_55_9 = 9;
  localparam control_matmul_55_10 = 10;
  localparam control_matmul_55_11 = 11;
  localparam control_matmul_55_12 = 12;
  localparam control_matmul_55_13 = 13;
  localparam control_matmul_55_14 = 14;
  localparam control_matmul_55_15 = 15;
  localparam control_matmul_55_16 = 16;
  localparam control_matmul_55_17 = 17;
  localparam control_matmul_55_18 = 18;
  localparam control_matmul_55_19 = 19;
  localparam control_matmul_55_20 = 20;
  localparam control_matmul_55_21 = 21;
  localparam control_matmul_55_22 = 22;
  localparam control_matmul_55_23 = 23;
  localparam control_matmul_55_24 = 24;
  localparam control_matmul_55_25 = 25;
  localparam control_matmul_55_26 = 26;
  localparam control_matmul_55_27 = 27;
  localparam control_matmul_55_28 = 28;

  always @(posedge CLK) begin
    if(RST) begin
      control_matmul_55 <= control_matmul_55_init;
      _control_matmul_55_called <= 0;
      matmul_55_filter_base_offset <= 0;
      matmul_55_filter_page_comp_offset <= 0;
      matmul_55_filter_page_dma_offset <= 0;
      matmul_55_act_base_offset_row <= 0;
      matmul_55_act_base_offset_bat <= 0;
      matmul_55_dma_flag_0 <= 0;
      matmul_55_act_page_comp_offset_0 <= 0;
      matmul_55_act_page_dma_offset_0 <= 0;
      matmul_55_out_base_offset_val <= 0;
      matmul_55_out_base_offset_col <= 0;
      matmul_55_out_base_offset_row <= 0;
      matmul_55_out_base_offset_bat <= 0;
      matmul_55_out_base_offset_och <= 0;
      matmul_55_out_page <= 0;
      matmul_55_out_page_comp_offset <= 0;
      matmul_55_out_page_dma_offset <= 0;
      matmul_55_out_laddr_offset <= 0;
      matmul_55_sync_out_count <= 0;
      matmul_55_write_count <= 0;
      matmul_55_next_out_write_size <= 0;
      matmul_55_row_count <= 0;
      matmul_55_bat_count <= 0;
      matmul_55_och_count <= 0;
      matmul_55_row_select <= 0;
      matmul_55_prev_row_count <= 0;
      matmul_55_prev_bat_count <= 0;
      matmul_55_prev_och_count <= 0;
      matmul_55_prev_row_select <= 0;
      matmul_55_out_col_count <= 0;
      matmul_55_out_row_count <= 0;
      matmul_55_out_ram_select <= 0;
      matmul_55_skip_read_filter <= 0;
      matmul_55_skip_read_act <= 0;
      matmul_55_skip_comp <= 0;
      matmul_55_skip_write_out <= 1;
    end else begin
      case(control_matmul_55)
        control_matmul_55_init: begin
          if(main_fsm == 134) begin
            _control_matmul_55_called <= 1;
          end 
          if(main_fsm == 144) begin
            _control_matmul_55_called <= 1;
          end 
          if(main_fsm == 154) begin
            _control_matmul_55_called <= 1;
          end 
          if(main_fsm == 134) begin
            control_matmul_55 <= control_matmul_55_1;
          end 
          if(main_fsm == 144) begin
            control_matmul_55 <= control_matmul_55_1;
          end 
          if(main_fsm == 154) begin
            control_matmul_55 <= control_matmul_55_1;
          end 
        end
        control_matmul_55_1: begin
          control_matmul_55 <= control_matmul_55_2;
        end
        control_matmul_55_2: begin
          matmul_55_filter_base_offset <= 0;
          matmul_55_filter_page_comp_offset <= 0;
          matmul_55_filter_page_dma_offset <= 0;
          matmul_55_act_base_offset_row <= 0;
          matmul_55_act_base_offset_bat <= 0;
          matmul_55_dma_flag_0 <= 1;
          matmul_55_act_page_comp_offset_0 <= 0;
          matmul_55_act_page_dma_offset_0 <= 0;
          matmul_55_out_base_offset_val <= 0;
          matmul_55_out_base_offset_col <= 0;
          matmul_55_out_base_offset_row <= 0;
          matmul_55_out_base_offset_bat <= 0;
          matmul_55_out_base_offset_och <= 0;
          matmul_55_out_page <= 0;
          matmul_55_out_page_comp_offset <= 0;
          matmul_55_out_page_dma_offset <= 0;
          matmul_55_out_laddr_offset <= 0;
          matmul_55_sync_out_count <= 0;
          matmul_55_write_count <= 0;
          matmul_55_next_out_write_size <= (cparam_matmul_55_max_och_count == 0)? cparam_matmul_55_out_write_size_res : cparam_matmul_55_out_write_size;
          matmul_55_row_count <= 0;
          matmul_55_bat_count <= 0;
          matmul_55_och_count <= 0;
          matmul_55_row_select <= 0;
          matmul_55_prev_row_count <= 0;
          matmul_55_prev_bat_count <= 0;
          matmul_55_prev_och_count <= 0;
          matmul_55_prev_row_select <= 0;
          matmul_55_out_col_count <= 0;
          matmul_55_out_row_count <= 0;
          matmul_55_out_ram_select <= 0;
          matmul_55_skip_read_filter <= 0;
          matmul_55_skip_read_act <= 0;
          matmul_55_skip_comp <= 0;
          matmul_55_skip_write_out <= 1;
          if(_maxi_read_req_idle) begin
            control_matmul_55 <= control_matmul_55_3;
          end 
        end
        control_matmul_55_3: begin
          if(_maxi_read_idle) begin
            control_matmul_55 <= control_matmul_55_4;
          end 
        end
        control_matmul_55_4: begin
          if(_maxi_read_req_idle) begin
            control_matmul_55 <= control_matmul_55_5;
          end 
        end
        control_matmul_55_5: begin
          if(_maxi_read_idle) begin
            control_matmul_55 <= control_matmul_55_6;
          end 
        end
        control_matmul_55_6: begin
          if(cparam_matmul_55_data_stationary == 0) begin
            control_matmul_55 <= control_matmul_55_7;
          end 
          if(cparam_matmul_55_data_stationary == 1) begin
            control_matmul_55 <= control_matmul_55_12;
          end 
        end
        control_matmul_55_7: begin
          control_matmul_55 <= control_matmul_55_8;
          if(matmul_55_skip_read_filter) begin
            control_matmul_55 <= control_matmul_55_11;
          end 
        end
        control_matmul_55_8: begin
          if(_maxi_read_req_idle) begin
            control_matmul_55 <= control_matmul_55_9;
          end 
        end
        control_matmul_55_9: begin
          if(_maxi_read_idle) begin
            control_matmul_55 <= control_matmul_55_10;
          end 
        end
        control_matmul_55_10: begin
          control_matmul_55 <= control_matmul_55_11;
        end
        control_matmul_55_11: begin
          if(cparam_matmul_55_data_stationary == 0) begin
            control_matmul_55 <= control_matmul_55_12;
          end 
          if(cparam_matmul_55_data_stationary == 1) begin
            control_matmul_55 <= control_matmul_55_18;
          end 
        end
        control_matmul_55_12: begin
          control_matmul_55 <= control_matmul_55_13;
          if(matmul_55_skip_read_act) begin
            control_matmul_55 <= control_matmul_55_17;
          end 
        end
        control_matmul_55_13: begin
          control_matmul_55 <= control_matmul_55_14;
          if(matmul_55_mux_dma_pad_mask_0 || !matmul_55_mux_dma_flag_0) begin
            control_matmul_55 <= control_matmul_55_16;
          end 
        end
        control_matmul_55_14: begin
          if(_maxi_read_req_idle) begin
            control_matmul_55 <= control_matmul_55_15;
          end 
        end
        control_matmul_55_15: begin
          if(_maxi_read_idle) begin
            control_matmul_55 <= control_matmul_55_16;
          end 
        end
        control_matmul_55_16: begin
          control_matmul_55 <= control_matmul_55_17;
        end
        control_matmul_55_17: begin
          if(cparam_matmul_55_data_stationary == 0) begin
            control_matmul_55 <= control_matmul_55_18;
          end 
          if(cparam_matmul_55_data_stationary == 1) begin
            control_matmul_55 <= control_matmul_55_7;
          end 
        end
        control_matmul_55_18: begin
          if(_maxi_write_idle) begin
            control_matmul_55 <= control_matmul_55_19;
          end 
        end
        control_matmul_55_19: begin
          if(matmul_55_comp_fsm == 0) begin
            control_matmul_55 <= control_matmul_55_20;
          end 
        end
        control_matmul_55_20: begin
          control_matmul_55 <= control_matmul_55_21;
          if(matmul_55_skip_write_out) begin
            control_matmul_55 <= control_matmul_55_26;
          end 
          if((cparam_matmul_55_data_stationary == 1) && (matmul_55_prev_och_count < cparam_matmul_55_max_och_count)) begin
            control_matmul_55 <= control_matmul_55_26;
          end 
        end
        control_matmul_55_21: begin
          if(matmul_55_sync_comp_count >= matmul_55_sync_out_count + cparam_matmul_55_inc_sync_out) begin
            control_matmul_55 <= control_matmul_55_22;
          end 
        end
        control_matmul_55_22: begin
          if(!matmul_55_dma_out_mask_0) begin
            control_matmul_55 <= control_matmul_55_23;
          end 
          if(matmul_55_dma_out_mask_0) begin
            control_matmul_55 <= control_matmul_55_24;
          end 
        end
        control_matmul_55_23: begin
          if(_maxi_write_req_idle) begin
            control_matmul_55 <= control_matmul_55_24;
          end 
        end
        control_matmul_55_24: begin
          control_matmul_55 <= control_matmul_55_25;
        end
        control_matmul_55_25: begin
          matmul_55_write_count <= matmul_55_write_count + 1;
          if(matmul_55_out_ram_select == 0) begin
            matmul_55_out_laddr_offset <= matmul_55_out_laddr_offset + matmul_55_next_out_write_size;
          end 
          if((cparam_matmul_55_data_stationary == 0) && !cparam_matmul_55_keep_filter) begin
            matmul_55_out_base_offset_col <= matmul_55_out_base_offset_col + cparam_matmul_55_out_col_step;
            matmul_55_out_col_count <= matmul_55_out_col_count + 1;
          end 
          matmul_55_out_ram_select <= matmul_55_out_ram_select + 1;
          if(matmul_55_out_ram_select == 0) begin
            matmul_55_out_ram_select <= 0;
          end 
          matmul_55_sync_out_count <= matmul_55_sync_out_count + cparam_matmul_55_inc_sync_out;
          if((cparam_matmul_55_data_stationary == 0) && !cparam_matmul_55_keep_filter && (matmul_55_write_count >= cparam_matmul_55_out_num_col - 1) || (cparam_matmul_55_data_stationary == 0) && cparam_matmul_55_keep_filter || (cparam_matmul_55_data_stationary == 1)) begin
            matmul_55_sync_out_count <= matmul_55_sync_out_count + (cparam_matmul_55_inc_sync_out + cparam_matmul_55_inc_sync_out_res);
          end 
          if((cparam_matmul_55_data_stationary == 0) && !cparam_matmul_55_keep_filter) begin
            control_matmul_55 <= control_matmul_55_20;
          end 
          if((cparam_matmul_55_data_stationary == 0) && !cparam_matmul_55_keep_filter && (matmul_55_write_count >= cparam_matmul_55_out_num_col - 1) || (cparam_matmul_55_data_stationary == 0) && cparam_matmul_55_keep_filter || (cparam_matmul_55_data_stationary == 1)) begin
            control_matmul_55 <= control_matmul_55_26;
          end 
        end
        control_matmul_55_26: begin
          if(matmul_55_update_filter) begin
            matmul_55_filter_base_offset <= matmul_55_filter_base_offset + cparam_matmul_55_filter_base_step;
          end 
          if((cparam_matmul_55_data_stationary == 1) && (matmul_55_och_count >= cparam_matmul_55_max_och_count)) begin
            matmul_55_filter_base_offset <= 0;
          end 
          if(matmul_55_update_filter) begin
            matmul_55_och_count <= matmul_55_och_count + cparam_matmul_55_och_count_step;
          end 
          if((cparam_matmul_55_data_stationary == 1) && (matmul_55_och_count >= cparam_matmul_55_max_och_count)) begin
            matmul_55_och_count <= 0;
          end 
          if(matmul_55_update_filter) begin
            matmul_55_filter_page_comp_offset <= matmul_55_filter_page_comp_offset + cparam_matmul_55_filter_read_step;
            matmul_55_filter_page_dma_offset <= matmul_55_filter_page_dma_offset + cparam_matmul_55_filter_read_step;
          end 
          if(matmul_55_update_filter && (matmul_55_filter_page_comp_offset + cparam_matmul_55_filter_read_step + cparam_matmul_55_filter_read_step > 262144)) begin
            matmul_55_filter_page_comp_offset <= 0;
            matmul_55_filter_page_dma_offset <= 0;
          end 
          if(matmul_55_update_act) begin
            matmul_55_act_base_offset_row <= matmul_55_act_base_offset_row + cparam_matmul_55_act_row_step;
          end 
          if(matmul_55_update_act && (matmul_55_row_count >= cparam_matmul_55_max_row_count)) begin
            matmul_55_act_base_offset_row <= 0;
            matmul_55_act_base_offset_bat <= matmul_55_act_base_offset_bat + cparam_matmul_55_act_bat_step;
          end 
          if(matmul_55_update_act && (matmul_55_row_count >= cparam_matmul_55_max_row_count) && (matmul_55_bat_count >= cparam_matmul_55_max_bat_count)) begin
            matmul_55_act_base_offset_bat <= 0;
          end 
          if(!matmul_55_update_act) begin
            matmul_55_dma_flag_0 <= 0;
          end 
          if(matmul_55_update_act) begin
            matmul_55_dma_flag_0 <= cparam_matmul_55_dma_flag_conds_0;
          end 
          if(matmul_55_update_act && (matmul_55_row_count >= cparam_matmul_55_max_row_count)) begin
            matmul_55_dma_flag_0 <= 1;
          end 
          if(matmul_55_update_act) begin
            matmul_55_row_count <= matmul_55_row_count + cparam_matmul_55_stride_row_par_row;
          end 
          if(matmul_55_update_act && (matmul_55_row_count >= cparam_matmul_55_max_row_count)) begin
            matmul_55_row_count <= 0;
            matmul_55_bat_count <= matmul_55_bat_count + 1;
          end 
          if(matmul_55_update_act && (matmul_55_row_count >= cparam_matmul_55_max_row_count) && (matmul_55_bat_count >= cparam_matmul_55_max_bat_count)) begin
            matmul_55_bat_count <= 0;
          end 
          if(matmul_55_update_act && (cparam_matmul_55_stride_row_par_row < 1)) begin
            matmul_55_row_select <= matmul_55_row_select + cparam_matmul_55_stride_row_par_row;
            matmul_55_prev_row_select <= matmul_55_row_select;
          end 
          if(matmul_55_update_act && (cparam_matmul_55_stride_row_par_row < 1) && (matmul_55_row_select + cparam_matmul_55_stride_row_par_row >= 1)) begin
            matmul_55_row_select <= matmul_55_row_select - (1 - cparam_matmul_55_stride_row_par_row);
            matmul_55_prev_row_select <= matmul_55_row_select;
          end 
          if(matmul_55_update_act && !(cparam_matmul_55_stride_row_par_row < 1)) begin
            matmul_55_row_select <= 0;
            matmul_55_prev_row_select <= 0;
          end 
          if(matmul_55_update_act && (matmul_55_row_count >= cparam_matmul_55_max_row_count)) begin
            matmul_55_row_select <= 0;
            matmul_55_prev_row_select <= 0;
          end 
          if(matmul_55_update_act && matmul_55_mux_next_dma_flag_0) begin
            matmul_55_act_page_comp_offset_0 <= matmul_55_act_page_comp_offset_0 + cparam_matmul_55_act_read_step;
            matmul_55_act_page_dma_offset_0 <= matmul_55_act_page_dma_offset_0 + cparam_matmul_55_act_read_step;
          end 
          if(matmul_55_update_act && matmul_55_mux_next_dma_flag_0 && (matmul_55_act_page_comp_offset_0 + cparam_matmul_55_act_read_step + cparam_matmul_55_act_read_step > 32768)) begin
            matmul_55_act_page_comp_offset_0 <= 0;
            matmul_55_act_page_dma_offset_0 <= 0;
          end 
          if((cparam_matmul_55_data_stationary == 0) && (matmul_55_row_count >= cparam_matmul_55_max_row_count) && (matmul_55_bat_count >= cparam_matmul_55_max_bat_count) && cparam_matmul_55_keep_input) begin
            matmul_55_act_page_comp_offset_0 <= 0;
            matmul_55_act_page_dma_offset_0 <= 0;
          end 
          matmul_55_next_out_write_size <= (matmul_55_och_count >= cparam_matmul_55_max_och_count)? cparam_matmul_55_out_write_size_res : cparam_matmul_55_out_write_size;
          if(!matmul_55_skip_write_out) begin
            matmul_55_write_count <= 0;
            matmul_55_out_laddr_offset <= 0;
            matmul_55_out_ram_select <= 0;
          end 
          if((cparam_matmul_55_data_stationary == 0) && !matmul_55_skip_write_out) begin
            matmul_55_out_base_offset_col <= 0;
            matmul_55_out_base_offset_row <= matmul_55_out_base_offset_row + cparam_matmul_55_out_row_step;
            matmul_55_out_col_count <= 0;
            matmul_55_out_row_count <= matmul_55_out_row_count + 1;
          end 
          if((cparam_matmul_55_data_stationary == 0) && !matmul_55_skip_write_out && (matmul_55_prev_row_count >= cparam_matmul_55_max_row_count)) begin
            matmul_55_out_base_offset_row <= 0;
            matmul_55_out_base_offset_bat <= matmul_55_out_base_offset_bat + cparam_matmul_55_out_bat_step;
            matmul_55_out_row_count <= 0;
          end 
          if((cparam_matmul_55_data_stationary == 0) && !matmul_55_skip_write_out && (matmul_55_prev_row_count >= cparam_matmul_55_max_row_count) && (matmul_55_prev_bat_count >= cparam_matmul_55_max_bat_count)) begin
            matmul_55_out_base_offset_bat <= 0;
            matmul_55_out_base_offset_och <= matmul_55_out_base_offset_och + cparam_matmul_55_out_och_step;
          end 
          if((cparam_matmul_55_data_stationary == 1) && (matmul_55_prev_och_count >= cparam_matmul_55_max_och_count) && !matmul_55_skip_write_out) begin
            matmul_55_out_base_offset_row <= matmul_55_out_base_offset_row + cparam_matmul_55_out_row_step;
          end 
          if((cparam_matmul_55_data_stationary == 0) && !matmul_55_out_page) begin
            matmul_55_out_page_comp_offset <= 1024;
            matmul_55_out_page_dma_offset <= 0;
            matmul_55_out_page <= 1;
          end 
          if((cparam_matmul_55_data_stationary == 0) && matmul_55_out_page) begin
            matmul_55_out_page_comp_offset <= 0;
            matmul_55_out_page_dma_offset <= 1024;
            matmul_55_out_page <= 0;
          end 
          if((cparam_matmul_55_data_stationary == 1) && (matmul_55_och_count >= cparam_matmul_55_max_och_count) && !matmul_55_out_page) begin
            matmul_55_out_page_comp_offset <= 1024;
            matmul_55_out_page_dma_offset <= 0;
            matmul_55_out_page <= 1;
          end 
          if((cparam_matmul_55_data_stationary == 1) && (matmul_55_och_count >= cparam_matmul_55_max_och_count) && matmul_55_out_page) begin
            matmul_55_out_page_comp_offset <= 0;
            matmul_55_out_page_dma_offset <= 1024;
            matmul_55_out_page <= 0;
          end 
          matmul_55_prev_row_count <= matmul_55_row_count;
          matmul_55_prev_bat_count <= matmul_55_bat_count;
          matmul_55_prev_och_count <= matmul_55_och_count;
          if((matmul_55_row_count >= cparam_matmul_55_max_row_count) && (matmul_55_bat_count >= cparam_matmul_55_max_bat_count) && (matmul_55_och_count >= cparam_matmul_55_max_och_count)) begin
            matmul_55_skip_read_filter <= 1;
          end 
          if((cparam_matmul_55_data_stationary == 1) && cparam_matmul_55_keep_filter) begin
            matmul_55_skip_read_filter <= 1;
          end 
          if((matmul_55_row_count >= cparam_matmul_55_max_row_count) && (matmul_55_bat_count >= cparam_matmul_55_max_bat_count) && (matmul_55_och_count >= cparam_matmul_55_max_och_count)) begin
            matmul_55_skip_read_act <= 1;
          end 
          if((cparam_matmul_55_data_stationary == 0) && (matmul_55_row_count >= cparam_matmul_55_max_row_count) && (matmul_55_bat_count >= cparam_matmul_55_max_bat_count) && cparam_matmul_55_keep_input) begin
            matmul_55_skip_read_act <= 1;
          end 
          if((matmul_55_row_count >= cparam_matmul_55_max_row_count) && (matmul_55_bat_count >= cparam_matmul_55_max_bat_count) && (matmul_55_och_count >= cparam_matmul_55_max_och_count)) begin
            matmul_55_skip_comp <= 1;
          end 
          if(matmul_55_skip_write_out && (matmul_55_prev_row_count == 0) && (matmul_55_prev_bat_count == 0) && (matmul_55_prev_och_count == 0)) begin
            matmul_55_skip_write_out <= 0;
          end 
          if(cparam_matmul_55_data_stationary == 0) begin
            control_matmul_55 <= control_matmul_55_12;
          end 
          if((cparam_matmul_55_data_stationary == 0) && (matmul_55_row_count >= cparam_matmul_55_max_row_count) && (matmul_55_bat_count >= cparam_matmul_55_max_bat_count)) begin
            control_matmul_55 <= control_matmul_55_7;
          end 
          if(cparam_matmul_55_data_stationary == 1) begin
            control_matmul_55 <= control_matmul_55_7;
          end 
          if((cparam_matmul_55_data_stationary == 1) && (matmul_55_och_count >= cparam_matmul_55_max_och_count)) begin
            control_matmul_55 <= control_matmul_55_12;
          end 
          if(!matmul_55_skip_write_out && (matmul_55_prev_och_count >= cparam_matmul_55_max_och_count) && (matmul_55_prev_row_count >= cparam_matmul_55_max_row_count) && (matmul_55_prev_bat_count >= cparam_matmul_55_max_bat_count)) begin
            control_matmul_55 <= control_matmul_55_27;
          end 
        end
        control_matmul_55_27: begin
          if(_maxi_write_idle && !_maxi_has_outstanding_write) begin
            control_matmul_55 <= control_matmul_55_28;
          end 
        end
        control_matmul_55_28: begin
          if(main_fsm == 137) begin
            _control_matmul_55_called <= 0;
          end 
          if(main_fsm == 147) begin
            _control_matmul_55_called <= 0;
          end 
          if(main_fsm == 157) begin
            _control_matmul_55_called <= 0;
          end 
          if(main_fsm == 137) begin
            control_matmul_55 <= control_matmul_55_init;
          end 
          if(main_fsm == 147) begin
            control_matmul_55 <= control_matmul_55_init;
          end 
          if(main_fsm == 157) begin
            control_matmul_55 <= control_matmul_55_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_29_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_29 <= write_burst_packed_fsm_29_init;
      write_burst_packed_addr_1644 <= 0;
      write_burst_packed_stride_1645 <= 0;
      write_burst_packed_length_1646 <= 0;
      write_burst_packed_done_1647 <= 0;
    end else begin
      case(write_burst_packed_fsm_29)
        write_burst_packed_fsm_29_init: begin
          write_burst_packed_addr_1644 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_1645 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_1646 <= _maxi_read_local_size_buf;
          write_burst_packed_done_1647 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 9) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_29 <= write_burst_packed_fsm_29_1;
          end 
        end
        write_burst_packed_fsm_29_1: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_packed_addr_1644 <= write_burst_packed_addr_1644 + write_burst_packed_stride_1645;
            write_burst_packed_length_1646 <= write_burst_packed_length_1646 - 1;
            write_burst_packed_done_1647 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_packed_length_1646 <= 1)) begin
            write_burst_packed_done_1647 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_packed_done_1647 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_packed_length_1646 <= 1)) begin
            write_burst_packed_fsm_29 <= write_burst_packed_fsm_29_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_packed_fsm_29 <= write_burst_packed_fsm_29_init;
          end 
          if(0) begin
            write_burst_packed_fsm_29 <= write_burst_packed_fsm_29_init;
          end 
        end
      endcase
    end
  end

  localparam matmul_55_comp_fsm_1 = 1;
  localparam matmul_55_comp_fsm_2 = 2;
  localparam matmul_55_comp_fsm_3 = 3;
  localparam matmul_55_comp_fsm_4 = 4;
  localparam matmul_55_comp_fsm_5 = 5;
  localparam matmul_55_comp_fsm_6 = 6;

  always @(posedge CLK) begin
    if(RST) begin
      matmul_55_comp_fsm <= matmul_55_comp_fsm_init;
      matmul_55_stream_act_local_0 <= 0;
      matmul_55_stream_out_local_col <= 0;
      matmul_55_stream_out_local_val <= 0;
      matmul_55_col_count <= 0;
      matmul_55_col_select <= 0;
      matmul_55_filter_page_comp_offset_buf <= 0;
      matmul_55_act_page_comp_offset_buf_0 <= 0;
      matmul_55_out_page_comp_offset_buf <= 0;
      matmul_55_row_count_buf <= 0;
      matmul_55_row_select_buf <= 0;
      matmul_55_och_count_buf <= 0;
      matmul_55_next_stream_num_ops <= 0;
      matmul_55_stream_pad_masks <= 0;
      matmul_55_sync_comp_count <= 0;
    end else begin
      if(_stream_matmul_55_sink_stop) begin
        matmul_55_sync_comp_count <= matmul_55_sync_comp_count + 1;
      end 
      if(control_matmul_55 == 6) begin
        matmul_55_sync_comp_count <= 0;
      end 
      case(matmul_55_comp_fsm)
        matmul_55_comp_fsm_init: begin
          if((control_matmul_55 == 19) && !matmul_55_skip_comp) begin
            matmul_55_comp_fsm <= matmul_55_comp_fsm_1;
          end 
        end
        matmul_55_comp_fsm_1: begin
          matmul_55_stream_act_local_0 <= 0;
          if(cparam_matmul_55_stream_act_local_small_flags_0) begin
            matmul_55_stream_act_local_0 <= cparam_matmul_55_stream_act_local_small_offset;
          end 
          if(cparam_matmul_55_stream_act_local_large_flags_0) begin
            matmul_55_stream_act_local_0 <= cparam_matmul_55_stream_act_local_large_offset;
          end 
          matmul_55_stream_out_local_col <= 0;
          if((cparam_matmul_55_data_stationary == 1) && (matmul_55_och_count == 0)) begin
            matmul_55_stream_out_local_val <= 0;
          end 
          matmul_55_col_count <= 0;
          matmul_55_col_select <= cparam_matmul_55_col_select_initval;
          matmul_55_filter_page_comp_offset_buf <= matmul_55_filter_page_comp_offset;
          matmul_55_act_page_comp_offset_buf_0 <= matmul_55_act_page_comp_offset_0;
          matmul_55_out_page_comp_offset_buf <= matmul_55_out_page_comp_offset;
          matmul_55_row_count_buf <= matmul_55_row_count;
          matmul_55_row_select_buf <= matmul_55_row_select;
          matmul_55_och_count_buf <= matmul_55_och_count;
          matmul_55_next_stream_num_ops <= (matmul_55_och_count >= cparam_matmul_55_max_och_count)? cparam_matmul_55_stream_num_ops_res : cparam_matmul_55_stream_num_ops;
          matmul_55_comp_fsm <= matmul_55_comp_fsm_2;
        end
        matmul_55_comp_fsm_2: begin
          matmul_55_stream_pad_masks <= { matmul_55_stream_pad_mask_0_0 };
          matmul_55_comp_fsm <= matmul_55_comp_fsm_3;
        end
        matmul_55_comp_fsm_3: begin
          matmul_55_comp_fsm <= matmul_55_comp_fsm_4;
          matmul_55_comp_fsm <= matmul_55_comp_fsm_4;
          matmul_55_comp_fsm <= matmul_55_comp_fsm_4;
          matmul_55_comp_fsm <= matmul_55_comp_fsm_4;
          matmul_55_comp_fsm <= matmul_55_comp_fsm_4;
          matmul_55_comp_fsm <= matmul_55_comp_fsm_4;
          matmul_55_comp_fsm <= matmul_55_comp_fsm_4;
          matmul_55_comp_fsm <= matmul_55_comp_fsm_4;
          matmul_55_comp_fsm <= matmul_55_comp_fsm_4;
          matmul_55_comp_fsm <= matmul_55_comp_fsm_4;
          matmul_55_comp_fsm <= matmul_55_comp_fsm_4;
          matmul_55_comp_fsm <= matmul_55_comp_fsm_4;
          matmul_55_comp_fsm <= matmul_55_comp_fsm_4;
          matmul_55_comp_fsm <= matmul_55_comp_fsm_4;
          matmul_55_comp_fsm <= matmul_55_comp_fsm_4;
          matmul_55_comp_fsm <= matmul_55_comp_fsm_4;
          matmul_55_comp_fsm <= matmul_55_comp_fsm_4;
          matmul_55_comp_fsm <= matmul_55_comp_fsm_4;
          matmul_55_comp_fsm <= matmul_55_comp_fsm_4;
          matmul_55_comp_fsm <= matmul_55_comp_fsm_4;
          matmul_55_comp_fsm <= matmul_55_comp_fsm_4;
          if(_stream_matmul_55_stream_oready) begin
            matmul_55_comp_fsm <= matmul_55_comp_fsm_4;
          end 
          matmul_55_comp_fsm <= matmul_55_comp_fsm_4;
        end
        matmul_55_comp_fsm_4: begin
          if(!_stream_matmul_55_source_busy) begin
            matmul_55_comp_fsm <= matmul_55_comp_fsm_5;
          end 
        end
        matmul_55_comp_fsm_5: begin
          if(_stream_matmul_55_busy) begin
            matmul_55_comp_fsm <= matmul_55_comp_fsm_6;
          end 
        end
        matmul_55_comp_fsm_6: begin
          if(!((matmul_55_col_select == 0)? cparam_matmul_55_inc_act_laddr_conds_0 : 0)) begin
            matmul_55_stream_act_local_0 <= matmul_55_stream_act_local_0 + cparam_matmul_55_inc_act_laddr_small;
          end 
          if((matmul_55_col_select == 0)? cparam_matmul_55_inc_act_laddr_conds_0 : 0) begin
            matmul_55_stream_act_local_0 <= matmul_55_stream_act_local_0 + cparam_matmul_55_inc_act_laddr_large;
          end 
          if(matmul_55_col_count >= cparam_matmul_55_max_col_count) begin
            matmul_55_stream_act_local_0 <= 0;
          end 
          if((matmul_55_col_count >= cparam_matmul_55_max_col_count) && cparam_matmul_55_stream_act_local_small_flags_0) begin
            matmul_55_stream_act_local_0 <= cparam_matmul_55_stream_act_local_small_offset;
          end 
          if((matmul_55_col_count >= cparam_matmul_55_max_col_count) && cparam_matmul_55_stream_act_local_large_flags_0) begin
            matmul_55_stream_act_local_0 <= cparam_matmul_55_stream_act_local_large_offset;
          end 
          if(cparam_matmul_55_data_stationary == 0) begin
            matmul_55_stream_out_local_col <= matmul_55_stream_out_local_col + matmul_55_next_stream_num_ops;
          end 
          if((cparam_matmul_55_data_stationary == 0) && (matmul_55_col_count >= cparam_matmul_55_max_col_count)) begin
            matmul_55_stream_out_local_col <= 0;
          end 
          if(cparam_matmul_55_data_stationary == 1) begin
            matmul_55_stream_out_local_col <= matmul_55_stream_out_local_col + cparam_matmul_55_inc_out_laddr_col;
          end 
          if((cparam_matmul_55_data_stationary == 1) && (matmul_55_col_count >= cparam_matmul_55_max_col_count)) begin
            matmul_55_stream_out_local_val <= matmul_55_stream_out_local_val + matmul_55_next_stream_num_ops;
            matmul_55_stream_out_local_col <= 0;
          end 
          matmul_55_col_count <= matmul_55_col_count + cparam_matmul_55_stride_col_par_col;
          if(matmul_55_col_count >= cparam_matmul_55_max_col_count) begin
            matmul_55_col_count <= 0;
          end 
          matmul_55_col_select <= matmul_55_col_select + cparam_matmul_55_stride_col_mod_filter_num;
          if(matmul_55_col_select + cparam_matmul_55_stride_col_mod_filter_num >= 1) begin
            matmul_55_col_select <= matmul_55_col_select - cparam_matmul_55_filter_num_col_minus_stride_col_mod;
          end 
          if(matmul_55_col_count >= cparam_matmul_55_max_col_count) begin
            matmul_55_col_select <= cparam_matmul_55_col_select_initval;
          end 
          matmul_55_comp_fsm <= matmul_55_comp_fsm_2;
          if(matmul_55_col_count >= cparam_matmul_55_max_col_count) begin
            matmul_55_comp_fsm <= matmul_55_comp_fsm_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_matmul_55_source_7_source_pat_fsm_0_1 = 1;
  localparam _stream_matmul_55_source_7_source_pat_fsm_0_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_matmul_55_source_7_source_pat_fsm_0 <= _stream_matmul_55_source_7_source_pat_fsm_0_init;
    end else begin
      case(_stream_matmul_55_source_7_source_pat_fsm_0)
        _stream_matmul_55_source_7_source_pat_fsm_0_init: begin
          if(_stream_matmul_55_source_start && _stream_matmul_55_source_7_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
            _stream_matmul_55_source_7_source_pat_fsm_0 <= _stream_matmul_55_source_7_source_pat_fsm_0_1;
          end 
        end
        _stream_matmul_55_source_7_source_pat_fsm_0_1: begin
          if(_stream_matmul_55_source_stop && _stream_matmul_55_stream_oready) begin
            _stream_matmul_55_source_7_source_pat_fsm_0 <= _stream_matmul_55_source_7_source_pat_fsm_0_init;
          end 
          if((_source_stream_matmul_55_source_7_pat_count_0 == 0) && (_source_stream_matmul_55_source_7_pat_count_1 == 0) && (_source_stream_matmul_55_source_7_pat_count_2 == 0) && (_source_stream_matmul_55_source_7_pat_count_3 == 0) && _stream_matmul_55_stream_oready) begin
            _stream_matmul_55_source_7_source_pat_fsm_0 <= _stream_matmul_55_source_7_source_pat_fsm_0_2;
          end 
        end
        _stream_matmul_55_source_7_source_pat_fsm_0_2: begin
          if(_stream_matmul_55_stream_oready) begin
            _stream_matmul_55_source_7_source_pat_fsm_0 <= _stream_matmul_55_source_7_source_pat_fsm_0_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_matmul_55_source_9_source_pat_fsm_1_1 = 1;
  localparam _stream_matmul_55_source_9_source_pat_fsm_1_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_matmul_55_source_9_source_pat_fsm_1 <= _stream_matmul_55_source_9_source_pat_fsm_1_init;
    end else begin
      case(_stream_matmul_55_source_9_source_pat_fsm_1)
        _stream_matmul_55_source_9_source_pat_fsm_1_init: begin
          if(_stream_matmul_55_source_start && _stream_matmul_55_source_9_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
            _stream_matmul_55_source_9_source_pat_fsm_1 <= _stream_matmul_55_source_9_source_pat_fsm_1_1;
          end 
        end
        _stream_matmul_55_source_9_source_pat_fsm_1_1: begin
          if(_stream_matmul_55_source_stop && _stream_matmul_55_stream_oready) begin
            _stream_matmul_55_source_9_source_pat_fsm_1 <= _stream_matmul_55_source_9_source_pat_fsm_1_init;
          end 
          if((_source_stream_matmul_55_source_9_pat_count_0 == 0) && (_source_stream_matmul_55_source_9_pat_count_1 == 0) && (_source_stream_matmul_55_source_9_pat_count_2 == 0) && (_source_stream_matmul_55_source_9_pat_count_3 == 0) && _stream_matmul_55_stream_oready) begin
            _stream_matmul_55_source_9_source_pat_fsm_1 <= _stream_matmul_55_source_9_source_pat_fsm_1_2;
          end 
        end
        _stream_matmul_55_source_9_source_pat_fsm_1_2: begin
          if(_stream_matmul_55_stream_oready) begin
            _stream_matmul_55_source_9_source_pat_fsm_1 <= _stream_matmul_55_source_9_source_pat_fsm_1_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_1691 <= 0;
    end else begin
      if(_stream_matmul_55_stream_oready && _stream_matmul_55_source_20_source_ram_renable && (_stream_matmul_55_source_20_source_sel == 3)) begin
        _tmp_1691 <= read_rtl_bank_1690;
      end 
    end
  end

  localparam _stream_matmul_55_source_20_source_pat_fsm_2_1 = 1;
  localparam _stream_matmul_55_source_20_source_pat_fsm_2_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_matmul_55_source_20_source_pat_fsm_2 <= _stream_matmul_55_source_20_source_pat_fsm_2_init;
    end else begin
      case(_stream_matmul_55_source_20_source_pat_fsm_2)
        _stream_matmul_55_source_20_source_pat_fsm_2_init: begin
          if(_stream_matmul_55_source_start && _stream_matmul_55_source_20_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
            _stream_matmul_55_source_20_source_pat_fsm_2 <= _stream_matmul_55_source_20_source_pat_fsm_2_1;
          end 
        end
        _stream_matmul_55_source_20_source_pat_fsm_2_1: begin
          if(_stream_matmul_55_source_stop && _stream_matmul_55_stream_oready) begin
            _stream_matmul_55_source_20_source_pat_fsm_2 <= _stream_matmul_55_source_20_source_pat_fsm_2_init;
          end 
          if((_source_stream_matmul_55_source_20_pat_count_0 == 0) && (_source_stream_matmul_55_source_20_pat_count_1 == 0) && (_source_stream_matmul_55_source_20_pat_count_2 == 0) && (_source_stream_matmul_55_source_20_pat_count_3 == 0) && _stream_matmul_55_stream_oready) begin
            _stream_matmul_55_source_20_source_pat_fsm_2 <= _stream_matmul_55_source_20_source_pat_fsm_2_2;
          end 
        end
        _stream_matmul_55_source_20_source_pat_fsm_2_2: begin
          if(_stream_matmul_55_stream_oready) begin
            _stream_matmul_55_source_20_source_pat_fsm_2 <= _stream_matmul_55_source_20_source_pat_fsm_2_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_matmul_55_source_21_source_pat_fsm_3_1 = 1;
  localparam _stream_matmul_55_source_21_source_pat_fsm_3_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_matmul_55_source_21_source_pat_fsm_3 <= _stream_matmul_55_source_21_source_pat_fsm_3_init;
    end else begin
      case(_stream_matmul_55_source_21_source_pat_fsm_3)
        _stream_matmul_55_source_21_source_pat_fsm_3_init: begin
          if(_stream_matmul_55_source_start && _stream_matmul_55_source_21_source_mode & 5'b10 && _stream_matmul_55_stream_oready) begin
            _stream_matmul_55_source_21_source_pat_fsm_3 <= _stream_matmul_55_source_21_source_pat_fsm_3_1;
          end 
        end
        _stream_matmul_55_source_21_source_pat_fsm_3_1: begin
          if(_stream_matmul_55_source_stop && _stream_matmul_55_stream_oready) begin
            _stream_matmul_55_source_21_source_pat_fsm_3 <= _stream_matmul_55_source_21_source_pat_fsm_3_init;
          end 
          if((_source_stream_matmul_55_source_21_pat_count_0 == 0) && (_source_stream_matmul_55_source_21_pat_count_1 == 0) && (_source_stream_matmul_55_source_21_pat_count_2 == 0) && (_source_stream_matmul_55_source_21_pat_count_3 == 0) && _stream_matmul_55_stream_oready) begin
            _stream_matmul_55_source_21_source_pat_fsm_3 <= _stream_matmul_55_source_21_source_pat_fsm_3_2;
          end 
        end
        _stream_matmul_55_source_21_source_pat_fsm_3_2: begin
          if(_stream_matmul_55_stream_oready) begin
            _stream_matmul_55_source_21_source_pat_fsm_3 <= _stream_matmul_55_source_21_source_pat_fsm_3_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_matmul_55_sink_26_sink_fsm_4_1 = 1;
  localparam _stream_matmul_55_sink_26_sink_fsm_4_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_matmul_55_sink_26_sink_fsm_4 <= _stream_matmul_55_sink_26_sink_fsm_4_init;
    end else begin
      case(_stream_matmul_55_sink_26_sink_fsm_4)
        _stream_matmul_55_sink_26_sink_fsm_4_init: begin
          if(_stream_matmul_55_sink_start && _stream_matmul_55_sink_26_sink_mode & 5'b1 && _stream_matmul_55_stream_oready) begin
            _stream_matmul_55_sink_26_sink_fsm_4 <= _stream_matmul_55_sink_26_sink_fsm_4_1;
          end 
        end
        _stream_matmul_55_sink_26_sink_fsm_4_1: begin
          if(_stream_matmul_55_stream_oready) begin
            _stream_matmul_55_sink_26_sink_fsm_4 <= _stream_matmul_55_sink_26_sink_fsm_4_2;
          end 
        end
        _stream_matmul_55_sink_26_sink_fsm_4_2: begin
          if(stream_matmul_55_sink_27_data && (_stream_matmul_55_sink_26_sink_count == 1) && _stream_matmul_55_stream_oready) begin
            _stream_matmul_55_sink_26_sink_fsm_4 <= _stream_matmul_55_sink_26_sink_fsm_4_init;
          end 
          if(_stream_matmul_55_sink_stop && _stream_matmul_55_stream_oready) begin
            _stream_matmul_55_sink_26_sink_fsm_4 <= _stream_matmul_55_sink_26_sink_fsm_4_init;
          end 
        end
      endcase
    end
  end


endmodule



module _maxi_read_req_fifo
(
  input CLK,
  input RST,
  input _maxi_read_req_fifo_enq,
  input [137-1:0] _maxi_read_req_fifo_wdata,
  output _maxi_read_req_fifo_full,
  output _maxi_read_req_fifo_almost_full,
  input _maxi_read_req_fifo_deq,
  output [137-1:0] _maxi_read_req_fifo_rdata,
  output _maxi_read_req_fifo_empty,
  output _maxi_read_req_fifo_almost_empty
);

  reg [137-1:0] mem [0:8-1];
  reg [3-1:0] head;
  reg [3-1:0] tail;
  wire is_empty;
  wire is_almost_empty;
  wire is_full;
  wire is_almost_full;
  assign is_empty = head == tail;
  assign is_almost_empty = head == (tail + 1 & 7);
  assign is_full = (head + 1 & 7) == tail;
  assign is_almost_full = (head + 2 & 7) == tail;
  wire [137-1:0] rdata;
  assign _maxi_read_req_fifo_full = is_full;
  assign _maxi_read_req_fifo_almost_full = is_almost_full || is_full;
  assign _maxi_read_req_fifo_empty = is_empty;
  assign _maxi_read_req_fifo_almost_empty = is_almost_empty || is_empty;
  assign rdata = mem[tail];
  assign _maxi_read_req_fifo_rdata = rdata;

  always @(posedge CLK) begin
    if(RST) begin
      head <= 0;
      tail <= 0;
    end else begin
      if(_maxi_read_req_fifo_enq && !is_full) begin
        mem[head] <= _maxi_read_req_fifo_wdata;
        head <= head + 1;
      end 
      if(_maxi_read_req_fifo_deq && !is_empty) begin
        tail <= tail + 1;
      end 
    end
  end


endmodule



module _maxi_write_req_fifo
(
  input CLK,
  input RST,
  input _maxi_write_req_fifo_enq,
  input [137-1:0] _maxi_write_req_fifo_wdata,
  output _maxi_write_req_fifo_full,
  output _maxi_write_req_fifo_almost_full,
  input _maxi_write_req_fifo_deq,
  output [137-1:0] _maxi_write_req_fifo_rdata,
  output _maxi_write_req_fifo_empty,
  output _maxi_write_req_fifo_almost_empty
);

  reg [137-1:0] mem [0:8-1];
  reg [3-1:0] head;
  reg [3-1:0] tail;
  wire is_empty;
  wire is_almost_empty;
  wire is_full;
  wire is_almost_full;
  assign is_empty = head == tail;
  assign is_almost_empty = head == (tail + 1 & 7);
  assign is_full = (head + 1 & 7) == tail;
  assign is_almost_full = (head + 2 & 7) == tail;
  wire [137-1:0] rdata;
  assign _maxi_write_req_fifo_full = is_full;
  assign _maxi_write_req_fifo_almost_full = is_almost_full || is_full;
  assign _maxi_write_req_fifo_empty = is_empty;
  assign _maxi_write_req_fifo_almost_empty = is_almost_empty || is_empty;
  assign rdata = mem[tail];
  assign _maxi_write_req_fifo_rdata = rdata;

  always @(posedge CLK) begin
    if(RST) begin
      head <= 0;
      tail <= 0;
    end else begin
      if(_maxi_write_req_fifo_enq && !is_full) begin
        mem[head] <= _maxi_write_req_fifo_wdata;
        head <= head + 1;
      end 
      if(_maxi_write_req_fifo_deq && !is_empty) begin
        tail <= tail + 1;
      end 
    end
  end


endmodule



module ram_w8_l262144_id0_0
(
  input CLK,
  input [16-1:0] ram_w8_l262144_id0_0_0_addr,
  output [8-1:0] ram_w8_l262144_id0_0_0_rdata,
  input [8-1:0] ram_w8_l262144_id0_0_0_wdata,
  input ram_w8_l262144_id0_0_0_wenable,
  input ram_w8_l262144_id0_0_0_enable,
  input [16-1:0] ram_w8_l262144_id0_0_1_addr,
  output [8-1:0] ram_w8_l262144_id0_0_1_rdata,
  input [8-1:0] ram_w8_l262144_id0_0_1_wdata,
  input ram_w8_l262144_id0_0_1_wenable,
  input ram_w8_l262144_id0_0_1_enable
);

  reg [8-1:0] ram_w8_l262144_id0_0_0_rdata_out;
  assign ram_w8_l262144_id0_0_0_rdata = ram_w8_l262144_id0_0_0_rdata_out;
  reg [8-1:0] ram_w8_l262144_id0_0_1_rdata_out;
  assign ram_w8_l262144_id0_0_1_rdata = ram_w8_l262144_id0_0_1_rdata_out;
  reg [8-1:0] mem [0:65536-1];

  always @(posedge CLK) begin
    if(ram_w8_l262144_id0_0_0_enable) begin
      if(ram_w8_l262144_id0_0_0_wenable) begin
        mem[ram_w8_l262144_id0_0_0_addr] <= ram_w8_l262144_id0_0_0_wdata;
        ram_w8_l262144_id0_0_0_rdata_out <= ram_w8_l262144_id0_0_0_wdata;
      end else begin
        ram_w8_l262144_id0_0_0_rdata_out <= mem[ram_w8_l262144_id0_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l262144_id0_0_1_enable) begin
      if(ram_w8_l262144_id0_0_1_wenable) begin
        mem[ram_w8_l262144_id0_0_1_addr] <= ram_w8_l262144_id0_0_1_wdata;
        ram_w8_l262144_id0_0_1_rdata_out <= ram_w8_l262144_id0_0_1_wdata;
      end else begin
        ram_w8_l262144_id0_0_1_rdata_out <= mem[ram_w8_l262144_id0_0_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l262144_id0_1
(
  input CLK,
  input [16-1:0] ram_w8_l262144_id0_1_0_addr,
  output [8-1:0] ram_w8_l262144_id0_1_0_rdata,
  input [8-1:0] ram_w8_l262144_id0_1_0_wdata,
  input ram_w8_l262144_id0_1_0_wenable,
  input ram_w8_l262144_id0_1_0_enable,
  input [16-1:0] ram_w8_l262144_id0_1_1_addr,
  output [8-1:0] ram_w8_l262144_id0_1_1_rdata,
  input [8-1:0] ram_w8_l262144_id0_1_1_wdata,
  input ram_w8_l262144_id0_1_1_wenable,
  input ram_w8_l262144_id0_1_1_enable
);

  reg [8-1:0] ram_w8_l262144_id0_1_0_rdata_out;
  assign ram_w8_l262144_id0_1_0_rdata = ram_w8_l262144_id0_1_0_rdata_out;
  reg [8-1:0] ram_w8_l262144_id0_1_1_rdata_out;
  assign ram_w8_l262144_id0_1_1_rdata = ram_w8_l262144_id0_1_1_rdata_out;
  reg [8-1:0] mem [0:65536-1];

  always @(posedge CLK) begin
    if(ram_w8_l262144_id0_1_0_enable) begin
      if(ram_w8_l262144_id0_1_0_wenable) begin
        mem[ram_w8_l262144_id0_1_0_addr] <= ram_w8_l262144_id0_1_0_wdata;
        ram_w8_l262144_id0_1_0_rdata_out <= ram_w8_l262144_id0_1_0_wdata;
      end else begin
        ram_w8_l262144_id0_1_0_rdata_out <= mem[ram_w8_l262144_id0_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l262144_id0_1_1_enable) begin
      if(ram_w8_l262144_id0_1_1_wenable) begin
        mem[ram_w8_l262144_id0_1_1_addr] <= ram_w8_l262144_id0_1_1_wdata;
        ram_w8_l262144_id0_1_1_rdata_out <= ram_w8_l262144_id0_1_1_wdata;
      end else begin
        ram_w8_l262144_id0_1_1_rdata_out <= mem[ram_w8_l262144_id0_1_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l262144_id0_2
(
  input CLK,
  input [16-1:0] ram_w8_l262144_id0_2_0_addr,
  output [8-1:0] ram_w8_l262144_id0_2_0_rdata,
  input [8-1:0] ram_w8_l262144_id0_2_0_wdata,
  input ram_w8_l262144_id0_2_0_wenable,
  input ram_w8_l262144_id0_2_0_enable,
  input [16-1:0] ram_w8_l262144_id0_2_1_addr,
  output [8-1:0] ram_w8_l262144_id0_2_1_rdata,
  input [8-1:0] ram_w8_l262144_id0_2_1_wdata,
  input ram_w8_l262144_id0_2_1_wenable,
  input ram_w8_l262144_id0_2_1_enable
);

  reg [8-1:0] ram_w8_l262144_id0_2_0_rdata_out;
  assign ram_w8_l262144_id0_2_0_rdata = ram_w8_l262144_id0_2_0_rdata_out;
  reg [8-1:0] ram_w8_l262144_id0_2_1_rdata_out;
  assign ram_w8_l262144_id0_2_1_rdata = ram_w8_l262144_id0_2_1_rdata_out;
  reg [8-1:0] mem [0:65536-1];

  always @(posedge CLK) begin
    if(ram_w8_l262144_id0_2_0_enable) begin
      if(ram_w8_l262144_id0_2_0_wenable) begin
        mem[ram_w8_l262144_id0_2_0_addr] <= ram_w8_l262144_id0_2_0_wdata;
        ram_w8_l262144_id0_2_0_rdata_out <= ram_w8_l262144_id0_2_0_wdata;
      end else begin
        ram_w8_l262144_id0_2_0_rdata_out <= mem[ram_w8_l262144_id0_2_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l262144_id0_2_1_enable) begin
      if(ram_w8_l262144_id0_2_1_wenable) begin
        mem[ram_w8_l262144_id0_2_1_addr] <= ram_w8_l262144_id0_2_1_wdata;
        ram_w8_l262144_id0_2_1_rdata_out <= ram_w8_l262144_id0_2_1_wdata;
      end else begin
        ram_w8_l262144_id0_2_1_rdata_out <= mem[ram_w8_l262144_id0_2_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l262144_id0_3
(
  input CLK,
  input [16-1:0] ram_w8_l262144_id0_3_0_addr,
  output [8-1:0] ram_w8_l262144_id0_3_0_rdata,
  input [8-1:0] ram_w8_l262144_id0_3_0_wdata,
  input ram_w8_l262144_id0_3_0_wenable,
  input ram_w8_l262144_id0_3_0_enable,
  input [16-1:0] ram_w8_l262144_id0_3_1_addr,
  output [8-1:0] ram_w8_l262144_id0_3_1_rdata,
  input [8-1:0] ram_w8_l262144_id0_3_1_wdata,
  input ram_w8_l262144_id0_3_1_wenable,
  input ram_w8_l262144_id0_3_1_enable
);

  reg [8-1:0] ram_w8_l262144_id0_3_0_rdata_out;
  assign ram_w8_l262144_id0_3_0_rdata = ram_w8_l262144_id0_3_0_rdata_out;
  reg [8-1:0] ram_w8_l262144_id0_3_1_rdata_out;
  assign ram_w8_l262144_id0_3_1_rdata = ram_w8_l262144_id0_3_1_rdata_out;
  reg [8-1:0] mem [0:65536-1];

  always @(posedge CLK) begin
    if(ram_w8_l262144_id0_3_0_enable) begin
      if(ram_w8_l262144_id0_3_0_wenable) begin
        mem[ram_w8_l262144_id0_3_0_addr] <= ram_w8_l262144_id0_3_0_wdata;
        ram_w8_l262144_id0_3_0_rdata_out <= ram_w8_l262144_id0_3_0_wdata;
      end else begin
        ram_w8_l262144_id0_3_0_rdata_out <= mem[ram_w8_l262144_id0_3_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l262144_id0_3_1_enable) begin
      if(ram_w8_l262144_id0_3_1_wenable) begin
        mem[ram_w8_l262144_id0_3_1_addr] <= ram_w8_l262144_id0_3_1_wdata;
        ram_w8_l262144_id0_3_1_rdata_out <= ram_w8_l262144_id0_3_1_wdata;
      end else begin
        ram_w8_l262144_id0_3_1_rdata_out <= mem[ram_w8_l262144_id0_3_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l32768_id0_0
(
  input CLK,
  input [13-1:0] ram_w8_l32768_id0_0_0_addr,
  output [8-1:0] ram_w8_l32768_id0_0_0_rdata,
  input [8-1:0] ram_w8_l32768_id0_0_0_wdata,
  input ram_w8_l32768_id0_0_0_wenable,
  input ram_w8_l32768_id0_0_0_enable,
  input [13-1:0] ram_w8_l32768_id0_0_1_addr,
  output [8-1:0] ram_w8_l32768_id0_0_1_rdata,
  input [8-1:0] ram_w8_l32768_id0_0_1_wdata,
  input ram_w8_l32768_id0_0_1_wenable,
  input ram_w8_l32768_id0_0_1_enable
);

  reg [8-1:0] ram_w8_l32768_id0_0_0_rdata_out;
  assign ram_w8_l32768_id0_0_0_rdata = ram_w8_l32768_id0_0_0_rdata_out;
  reg [8-1:0] ram_w8_l32768_id0_0_1_rdata_out;
  assign ram_w8_l32768_id0_0_1_rdata = ram_w8_l32768_id0_0_1_rdata_out;
  reg [8-1:0] mem [0:8192-1];

  always @(posedge CLK) begin
    if(ram_w8_l32768_id0_0_0_enable) begin
      if(ram_w8_l32768_id0_0_0_wenable) begin
        mem[ram_w8_l32768_id0_0_0_addr] <= ram_w8_l32768_id0_0_0_wdata;
        ram_w8_l32768_id0_0_0_rdata_out <= ram_w8_l32768_id0_0_0_wdata;
      end else begin
        ram_w8_l32768_id0_0_0_rdata_out <= mem[ram_w8_l32768_id0_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l32768_id0_0_1_enable) begin
      if(ram_w8_l32768_id0_0_1_wenable) begin
        mem[ram_w8_l32768_id0_0_1_addr] <= ram_w8_l32768_id0_0_1_wdata;
        ram_w8_l32768_id0_0_1_rdata_out <= ram_w8_l32768_id0_0_1_wdata;
      end else begin
        ram_w8_l32768_id0_0_1_rdata_out <= mem[ram_w8_l32768_id0_0_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l32768_id0_1
(
  input CLK,
  input [13-1:0] ram_w8_l32768_id0_1_0_addr,
  output [8-1:0] ram_w8_l32768_id0_1_0_rdata,
  input [8-1:0] ram_w8_l32768_id0_1_0_wdata,
  input ram_w8_l32768_id0_1_0_wenable,
  input ram_w8_l32768_id0_1_0_enable,
  input [13-1:0] ram_w8_l32768_id0_1_1_addr,
  output [8-1:0] ram_w8_l32768_id0_1_1_rdata,
  input [8-1:0] ram_w8_l32768_id0_1_1_wdata,
  input ram_w8_l32768_id0_1_1_wenable,
  input ram_w8_l32768_id0_1_1_enable
);

  reg [8-1:0] ram_w8_l32768_id0_1_0_rdata_out;
  assign ram_w8_l32768_id0_1_0_rdata = ram_w8_l32768_id0_1_0_rdata_out;
  reg [8-1:0] ram_w8_l32768_id0_1_1_rdata_out;
  assign ram_w8_l32768_id0_1_1_rdata = ram_w8_l32768_id0_1_1_rdata_out;
  reg [8-1:0] mem [0:8192-1];

  always @(posedge CLK) begin
    if(ram_w8_l32768_id0_1_0_enable) begin
      if(ram_w8_l32768_id0_1_0_wenable) begin
        mem[ram_w8_l32768_id0_1_0_addr] <= ram_w8_l32768_id0_1_0_wdata;
        ram_w8_l32768_id0_1_0_rdata_out <= ram_w8_l32768_id0_1_0_wdata;
      end else begin
        ram_w8_l32768_id0_1_0_rdata_out <= mem[ram_w8_l32768_id0_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l32768_id0_1_1_enable) begin
      if(ram_w8_l32768_id0_1_1_wenable) begin
        mem[ram_w8_l32768_id0_1_1_addr] <= ram_w8_l32768_id0_1_1_wdata;
        ram_w8_l32768_id0_1_1_rdata_out <= ram_w8_l32768_id0_1_1_wdata;
      end else begin
        ram_w8_l32768_id0_1_1_rdata_out <= mem[ram_w8_l32768_id0_1_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l32768_id0_2
(
  input CLK,
  input [13-1:0] ram_w8_l32768_id0_2_0_addr,
  output [8-1:0] ram_w8_l32768_id0_2_0_rdata,
  input [8-1:0] ram_w8_l32768_id0_2_0_wdata,
  input ram_w8_l32768_id0_2_0_wenable,
  input ram_w8_l32768_id0_2_0_enable,
  input [13-1:0] ram_w8_l32768_id0_2_1_addr,
  output [8-1:0] ram_w8_l32768_id0_2_1_rdata,
  input [8-1:0] ram_w8_l32768_id0_2_1_wdata,
  input ram_w8_l32768_id0_2_1_wenable,
  input ram_w8_l32768_id0_2_1_enable
);

  reg [8-1:0] ram_w8_l32768_id0_2_0_rdata_out;
  assign ram_w8_l32768_id0_2_0_rdata = ram_w8_l32768_id0_2_0_rdata_out;
  reg [8-1:0] ram_w8_l32768_id0_2_1_rdata_out;
  assign ram_w8_l32768_id0_2_1_rdata = ram_w8_l32768_id0_2_1_rdata_out;
  reg [8-1:0] mem [0:8192-1];

  always @(posedge CLK) begin
    if(ram_w8_l32768_id0_2_0_enable) begin
      if(ram_w8_l32768_id0_2_0_wenable) begin
        mem[ram_w8_l32768_id0_2_0_addr] <= ram_w8_l32768_id0_2_0_wdata;
        ram_w8_l32768_id0_2_0_rdata_out <= ram_w8_l32768_id0_2_0_wdata;
      end else begin
        ram_w8_l32768_id0_2_0_rdata_out <= mem[ram_w8_l32768_id0_2_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l32768_id0_2_1_enable) begin
      if(ram_w8_l32768_id0_2_1_wenable) begin
        mem[ram_w8_l32768_id0_2_1_addr] <= ram_w8_l32768_id0_2_1_wdata;
        ram_w8_l32768_id0_2_1_rdata_out <= ram_w8_l32768_id0_2_1_wdata;
      end else begin
        ram_w8_l32768_id0_2_1_rdata_out <= mem[ram_w8_l32768_id0_2_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l32768_id0_3
(
  input CLK,
  input [13-1:0] ram_w8_l32768_id0_3_0_addr,
  output [8-1:0] ram_w8_l32768_id0_3_0_rdata,
  input [8-1:0] ram_w8_l32768_id0_3_0_wdata,
  input ram_w8_l32768_id0_3_0_wenable,
  input ram_w8_l32768_id0_3_0_enable,
  input [13-1:0] ram_w8_l32768_id0_3_1_addr,
  output [8-1:0] ram_w8_l32768_id0_3_1_rdata,
  input [8-1:0] ram_w8_l32768_id0_3_1_wdata,
  input ram_w8_l32768_id0_3_1_wenable,
  input ram_w8_l32768_id0_3_1_enable
);

  reg [8-1:0] ram_w8_l32768_id0_3_0_rdata_out;
  assign ram_w8_l32768_id0_3_0_rdata = ram_w8_l32768_id0_3_0_rdata_out;
  reg [8-1:0] ram_w8_l32768_id0_3_1_rdata_out;
  assign ram_w8_l32768_id0_3_1_rdata = ram_w8_l32768_id0_3_1_rdata_out;
  reg [8-1:0] mem [0:8192-1];

  always @(posedge CLK) begin
    if(ram_w8_l32768_id0_3_0_enable) begin
      if(ram_w8_l32768_id0_3_0_wenable) begin
        mem[ram_w8_l32768_id0_3_0_addr] <= ram_w8_l32768_id0_3_0_wdata;
        ram_w8_l32768_id0_3_0_rdata_out <= ram_w8_l32768_id0_3_0_wdata;
      end else begin
        ram_w8_l32768_id0_3_0_rdata_out <= mem[ram_w8_l32768_id0_3_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l32768_id0_3_1_enable) begin
      if(ram_w8_l32768_id0_3_1_wenable) begin
        mem[ram_w8_l32768_id0_3_1_addr] <= ram_w8_l32768_id0_3_1_wdata;
        ram_w8_l32768_id0_3_1_rdata_out <= ram_w8_l32768_id0_3_1_wdata;
      end else begin
        ram_w8_l32768_id0_3_1_rdata_out <= mem[ram_w8_l32768_id0_3_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l16384_id0_0
(
  input CLK,
  input [12-1:0] ram_w8_l16384_id0_0_0_addr,
  output [8-1:0] ram_w8_l16384_id0_0_0_rdata,
  input [8-1:0] ram_w8_l16384_id0_0_0_wdata,
  input ram_w8_l16384_id0_0_0_wenable,
  input ram_w8_l16384_id0_0_0_enable,
  input [12-1:0] ram_w8_l16384_id0_0_1_addr,
  output [8-1:0] ram_w8_l16384_id0_0_1_rdata,
  input [8-1:0] ram_w8_l16384_id0_0_1_wdata,
  input ram_w8_l16384_id0_0_1_wenable,
  input ram_w8_l16384_id0_0_1_enable
);

  reg [8-1:0] ram_w8_l16384_id0_0_0_rdata_out;
  assign ram_w8_l16384_id0_0_0_rdata = ram_w8_l16384_id0_0_0_rdata_out;
  reg [8-1:0] ram_w8_l16384_id0_0_1_rdata_out;
  assign ram_w8_l16384_id0_0_1_rdata = ram_w8_l16384_id0_0_1_rdata_out;
  reg [8-1:0] mem [0:4096-1];

  always @(posedge CLK) begin
    if(ram_w8_l16384_id0_0_0_enable) begin
      if(ram_w8_l16384_id0_0_0_wenable) begin
        mem[ram_w8_l16384_id0_0_0_addr] <= ram_w8_l16384_id0_0_0_wdata;
        ram_w8_l16384_id0_0_0_rdata_out <= ram_w8_l16384_id0_0_0_wdata;
      end else begin
        ram_w8_l16384_id0_0_0_rdata_out <= mem[ram_w8_l16384_id0_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l16384_id0_0_1_enable) begin
      if(ram_w8_l16384_id0_0_1_wenable) begin
        mem[ram_w8_l16384_id0_0_1_addr] <= ram_w8_l16384_id0_0_1_wdata;
        ram_w8_l16384_id0_0_1_rdata_out <= ram_w8_l16384_id0_0_1_wdata;
      end else begin
        ram_w8_l16384_id0_0_1_rdata_out <= mem[ram_w8_l16384_id0_0_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l16384_id0_1
(
  input CLK,
  input [12-1:0] ram_w8_l16384_id0_1_0_addr,
  output [8-1:0] ram_w8_l16384_id0_1_0_rdata,
  input [8-1:0] ram_w8_l16384_id0_1_0_wdata,
  input ram_w8_l16384_id0_1_0_wenable,
  input ram_w8_l16384_id0_1_0_enable,
  input [12-1:0] ram_w8_l16384_id0_1_1_addr,
  output [8-1:0] ram_w8_l16384_id0_1_1_rdata,
  input [8-1:0] ram_w8_l16384_id0_1_1_wdata,
  input ram_w8_l16384_id0_1_1_wenable,
  input ram_w8_l16384_id0_1_1_enable
);

  reg [8-1:0] ram_w8_l16384_id0_1_0_rdata_out;
  assign ram_w8_l16384_id0_1_0_rdata = ram_w8_l16384_id0_1_0_rdata_out;
  reg [8-1:0] ram_w8_l16384_id0_1_1_rdata_out;
  assign ram_w8_l16384_id0_1_1_rdata = ram_w8_l16384_id0_1_1_rdata_out;
  reg [8-1:0] mem [0:4096-1];

  always @(posedge CLK) begin
    if(ram_w8_l16384_id0_1_0_enable) begin
      if(ram_w8_l16384_id0_1_0_wenable) begin
        mem[ram_w8_l16384_id0_1_0_addr] <= ram_w8_l16384_id0_1_0_wdata;
        ram_w8_l16384_id0_1_0_rdata_out <= ram_w8_l16384_id0_1_0_wdata;
      end else begin
        ram_w8_l16384_id0_1_0_rdata_out <= mem[ram_w8_l16384_id0_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l16384_id0_1_1_enable) begin
      if(ram_w8_l16384_id0_1_1_wenable) begin
        mem[ram_w8_l16384_id0_1_1_addr] <= ram_w8_l16384_id0_1_1_wdata;
        ram_w8_l16384_id0_1_1_rdata_out <= ram_w8_l16384_id0_1_1_wdata;
      end else begin
        ram_w8_l16384_id0_1_1_rdata_out <= mem[ram_w8_l16384_id0_1_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l16384_id0_2
(
  input CLK,
  input [12-1:0] ram_w8_l16384_id0_2_0_addr,
  output [8-1:0] ram_w8_l16384_id0_2_0_rdata,
  input [8-1:0] ram_w8_l16384_id0_2_0_wdata,
  input ram_w8_l16384_id0_2_0_wenable,
  input ram_w8_l16384_id0_2_0_enable,
  input [12-1:0] ram_w8_l16384_id0_2_1_addr,
  output [8-1:0] ram_w8_l16384_id0_2_1_rdata,
  input [8-1:0] ram_w8_l16384_id0_2_1_wdata,
  input ram_w8_l16384_id0_2_1_wenable,
  input ram_w8_l16384_id0_2_1_enable
);

  reg [8-1:0] ram_w8_l16384_id0_2_0_rdata_out;
  assign ram_w8_l16384_id0_2_0_rdata = ram_w8_l16384_id0_2_0_rdata_out;
  reg [8-1:0] ram_w8_l16384_id0_2_1_rdata_out;
  assign ram_w8_l16384_id0_2_1_rdata = ram_w8_l16384_id0_2_1_rdata_out;
  reg [8-1:0] mem [0:4096-1];

  always @(posedge CLK) begin
    if(ram_w8_l16384_id0_2_0_enable) begin
      if(ram_w8_l16384_id0_2_0_wenable) begin
        mem[ram_w8_l16384_id0_2_0_addr] <= ram_w8_l16384_id0_2_0_wdata;
        ram_w8_l16384_id0_2_0_rdata_out <= ram_w8_l16384_id0_2_0_wdata;
      end else begin
        ram_w8_l16384_id0_2_0_rdata_out <= mem[ram_w8_l16384_id0_2_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l16384_id0_2_1_enable) begin
      if(ram_w8_l16384_id0_2_1_wenable) begin
        mem[ram_w8_l16384_id0_2_1_addr] <= ram_w8_l16384_id0_2_1_wdata;
        ram_w8_l16384_id0_2_1_rdata_out <= ram_w8_l16384_id0_2_1_wdata;
      end else begin
        ram_w8_l16384_id0_2_1_rdata_out <= mem[ram_w8_l16384_id0_2_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l16384_id0_3
(
  input CLK,
  input [12-1:0] ram_w8_l16384_id0_3_0_addr,
  output [8-1:0] ram_w8_l16384_id0_3_0_rdata,
  input [8-1:0] ram_w8_l16384_id0_3_0_wdata,
  input ram_w8_l16384_id0_3_0_wenable,
  input ram_w8_l16384_id0_3_0_enable,
  input [12-1:0] ram_w8_l16384_id0_3_1_addr,
  output [8-1:0] ram_w8_l16384_id0_3_1_rdata,
  input [8-1:0] ram_w8_l16384_id0_3_1_wdata,
  input ram_w8_l16384_id0_3_1_wenable,
  input ram_w8_l16384_id0_3_1_enable
);

  reg [8-1:0] ram_w8_l16384_id0_3_0_rdata_out;
  assign ram_w8_l16384_id0_3_0_rdata = ram_w8_l16384_id0_3_0_rdata_out;
  reg [8-1:0] ram_w8_l16384_id0_3_1_rdata_out;
  assign ram_w8_l16384_id0_3_1_rdata = ram_w8_l16384_id0_3_1_rdata_out;
  reg [8-1:0] mem [0:4096-1];

  always @(posedge CLK) begin
    if(ram_w8_l16384_id0_3_0_enable) begin
      if(ram_w8_l16384_id0_3_0_wenable) begin
        mem[ram_w8_l16384_id0_3_0_addr] <= ram_w8_l16384_id0_3_0_wdata;
        ram_w8_l16384_id0_3_0_rdata_out <= ram_w8_l16384_id0_3_0_wdata;
      end else begin
        ram_w8_l16384_id0_3_0_rdata_out <= mem[ram_w8_l16384_id0_3_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l16384_id0_3_1_enable) begin
      if(ram_w8_l16384_id0_3_1_wenable) begin
        mem[ram_w8_l16384_id0_3_1_addr] <= ram_w8_l16384_id0_3_1_wdata;
        ram_w8_l16384_id0_3_1_rdata_out <= ram_w8_l16384_id0_3_1_wdata;
      end else begin
        ram_w8_l16384_id0_3_1_rdata_out <= mem[ram_w8_l16384_id0_3_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l16384_id1_0
(
  input CLK,
  input [12-1:0] ram_w8_l16384_id1_0_0_addr,
  output [8-1:0] ram_w8_l16384_id1_0_0_rdata,
  input [8-1:0] ram_w8_l16384_id1_0_0_wdata,
  input ram_w8_l16384_id1_0_0_wenable,
  input ram_w8_l16384_id1_0_0_enable,
  input [12-1:0] ram_w8_l16384_id1_0_1_addr,
  output [8-1:0] ram_w8_l16384_id1_0_1_rdata,
  input [8-1:0] ram_w8_l16384_id1_0_1_wdata,
  input ram_w8_l16384_id1_0_1_wenable,
  input ram_w8_l16384_id1_0_1_enable
);

  reg [8-1:0] ram_w8_l16384_id1_0_0_rdata_out;
  assign ram_w8_l16384_id1_0_0_rdata = ram_w8_l16384_id1_0_0_rdata_out;
  reg [8-1:0] ram_w8_l16384_id1_0_1_rdata_out;
  assign ram_w8_l16384_id1_0_1_rdata = ram_w8_l16384_id1_0_1_rdata_out;
  reg [8-1:0] mem [0:4096-1];

  always @(posedge CLK) begin
    if(ram_w8_l16384_id1_0_0_enable) begin
      if(ram_w8_l16384_id1_0_0_wenable) begin
        mem[ram_w8_l16384_id1_0_0_addr] <= ram_w8_l16384_id1_0_0_wdata;
        ram_w8_l16384_id1_0_0_rdata_out <= ram_w8_l16384_id1_0_0_wdata;
      end else begin
        ram_w8_l16384_id1_0_0_rdata_out <= mem[ram_w8_l16384_id1_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l16384_id1_0_1_enable) begin
      if(ram_w8_l16384_id1_0_1_wenable) begin
        mem[ram_w8_l16384_id1_0_1_addr] <= ram_w8_l16384_id1_0_1_wdata;
        ram_w8_l16384_id1_0_1_rdata_out <= ram_w8_l16384_id1_0_1_wdata;
      end else begin
        ram_w8_l16384_id1_0_1_rdata_out <= mem[ram_w8_l16384_id1_0_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l16384_id1_1
(
  input CLK,
  input [12-1:0] ram_w8_l16384_id1_1_0_addr,
  output [8-1:0] ram_w8_l16384_id1_1_0_rdata,
  input [8-1:0] ram_w8_l16384_id1_1_0_wdata,
  input ram_w8_l16384_id1_1_0_wenable,
  input ram_w8_l16384_id1_1_0_enable,
  input [12-1:0] ram_w8_l16384_id1_1_1_addr,
  output [8-1:0] ram_w8_l16384_id1_1_1_rdata,
  input [8-1:0] ram_w8_l16384_id1_1_1_wdata,
  input ram_w8_l16384_id1_1_1_wenable,
  input ram_w8_l16384_id1_1_1_enable
);

  reg [8-1:0] ram_w8_l16384_id1_1_0_rdata_out;
  assign ram_w8_l16384_id1_1_0_rdata = ram_w8_l16384_id1_1_0_rdata_out;
  reg [8-1:0] ram_w8_l16384_id1_1_1_rdata_out;
  assign ram_w8_l16384_id1_1_1_rdata = ram_w8_l16384_id1_1_1_rdata_out;
  reg [8-1:0] mem [0:4096-1];

  always @(posedge CLK) begin
    if(ram_w8_l16384_id1_1_0_enable) begin
      if(ram_w8_l16384_id1_1_0_wenable) begin
        mem[ram_w8_l16384_id1_1_0_addr] <= ram_w8_l16384_id1_1_0_wdata;
        ram_w8_l16384_id1_1_0_rdata_out <= ram_w8_l16384_id1_1_0_wdata;
      end else begin
        ram_w8_l16384_id1_1_0_rdata_out <= mem[ram_w8_l16384_id1_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l16384_id1_1_1_enable) begin
      if(ram_w8_l16384_id1_1_1_wenable) begin
        mem[ram_w8_l16384_id1_1_1_addr] <= ram_w8_l16384_id1_1_1_wdata;
        ram_w8_l16384_id1_1_1_rdata_out <= ram_w8_l16384_id1_1_1_wdata;
      end else begin
        ram_w8_l16384_id1_1_1_rdata_out <= mem[ram_w8_l16384_id1_1_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l16384_id1_2
(
  input CLK,
  input [12-1:0] ram_w8_l16384_id1_2_0_addr,
  output [8-1:0] ram_w8_l16384_id1_2_0_rdata,
  input [8-1:0] ram_w8_l16384_id1_2_0_wdata,
  input ram_w8_l16384_id1_2_0_wenable,
  input ram_w8_l16384_id1_2_0_enable,
  input [12-1:0] ram_w8_l16384_id1_2_1_addr,
  output [8-1:0] ram_w8_l16384_id1_2_1_rdata,
  input [8-1:0] ram_w8_l16384_id1_2_1_wdata,
  input ram_w8_l16384_id1_2_1_wenable,
  input ram_w8_l16384_id1_2_1_enable
);

  reg [8-1:0] ram_w8_l16384_id1_2_0_rdata_out;
  assign ram_w8_l16384_id1_2_0_rdata = ram_w8_l16384_id1_2_0_rdata_out;
  reg [8-1:0] ram_w8_l16384_id1_2_1_rdata_out;
  assign ram_w8_l16384_id1_2_1_rdata = ram_w8_l16384_id1_2_1_rdata_out;
  reg [8-1:0] mem [0:4096-1];

  always @(posedge CLK) begin
    if(ram_w8_l16384_id1_2_0_enable) begin
      if(ram_w8_l16384_id1_2_0_wenable) begin
        mem[ram_w8_l16384_id1_2_0_addr] <= ram_w8_l16384_id1_2_0_wdata;
        ram_w8_l16384_id1_2_0_rdata_out <= ram_w8_l16384_id1_2_0_wdata;
      end else begin
        ram_w8_l16384_id1_2_0_rdata_out <= mem[ram_w8_l16384_id1_2_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l16384_id1_2_1_enable) begin
      if(ram_w8_l16384_id1_2_1_wenable) begin
        mem[ram_w8_l16384_id1_2_1_addr] <= ram_w8_l16384_id1_2_1_wdata;
        ram_w8_l16384_id1_2_1_rdata_out <= ram_w8_l16384_id1_2_1_wdata;
      end else begin
        ram_w8_l16384_id1_2_1_rdata_out <= mem[ram_w8_l16384_id1_2_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l16384_id1_3
(
  input CLK,
  input [12-1:0] ram_w8_l16384_id1_3_0_addr,
  output [8-1:0] ram_w8_l16384_id1_3_0_rdata,
  input [8-1:0] ram_w8_l16384_id1_3_0_wdata,
  input ram_w8_l16384_id1_3_0_wenable,
  input ram_w8_l16384_id1_3_0_enable,
  input [12-1:0] ram_w8_l16384_id1_3_1_addr,
  output [8-1:0] ram_w8_l16384_id1_3_1_rdata,
  input [8-1:0] ram_w8_l16384_id1_3_1_wdata,
  input ram_w8_l16384_id1_3_1_wenable,
  input ram_w8_l16384_id1_3_1_enable
);

  reg [8-1:0] ram_w8_l16384_id1_3_0_rdata_out;
  assign ram_w8_l16384_id1_3_0_rdata = ram_w8_l16384_id1_3_0_rdata_out;
  reg [8-1:0] ram_w8_l16384_id1_3_1_rdata_out;
  assign ram_w8_l16384_id1_3_1_rdata = ram_w8_l16384_id1_3_1_rdata_out;
  reg [8-1:0] mem [0:4096-1];

  always @(posedge CLK) begin
    if(ram_w8_l16384_id1_3_0_enable) begin
      if(ram_w8_l16384_id1_3_0_wenable) begin
        mem[ram_w8_l16384_id1_3_0_addr] <= ram_w8_l16384_id1_3_0_wdata;
        ram_w8_l16384_id1_3_0_rdata_out <= ram_w8_l16384_id1_3_0_wdata;
      end else begin
        ram_w8_l16384_id1_3_0_rdata_out <= mem[ram_w8_l16384_id1_3_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l16384_id1_3_1_enable) begin
      if(ram_w8_l16384_id1_3_1_wenable) begin
        mem[ram_w8_l16384_id1_3_1_addr] <= ram_w8_l16384_id1_3_1_wdata;
        ram_w8_l16384_id1_3_1_rdata_out <= ram_w8_l16384_id1_3_1_wdata;
      end else begin
        ram_w8_l16384_id1_3_1_rdata_out <= mem[ram_w8_l16384_id1_3_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l16384_id2_0
(
  input CLK,
  input [12-1:0] ram_w8_l16384_id2_0_0_addr,
  output [8-1:0] ram_w8_l16384_id2_0_0_rdata,
  input [8-1:0] ram_w8_l16384_id2_0_0_wdata,
  input ram_w8_l16384_id2_0_0_wenable,
  input ram_w8_l16384_id2_0_0_enable,
  input [12-1:0] ram_w8_l16384_id2_0_1_addr,
  output [8-1:0] ram_w8_l16384_id2_0_1_rdata,
  input [8-1:0] ram_w8_l16384_id2_0_1_wdata,
  input ram_w8_l16384_id2_0_1_wenable,
  input ram_w8_l16384_id2_0_1_enable
);

  reg [8-1:0] ram_w8_l16384_id2_0_0_rdata_out;
  assign ram_w8_l16384_id2_0_0_rdata = ram_w8_l16384_id2_0_0_rdata_out;
  reg [8-1:0] ram_w8_l16384_id2_0_1_rdata_out;
  assign ram_w8_l16384_id2_0_1_rdata = ram_w8_l16384_id2_0_1_rdata_out;
  reg [8-1:0] mem [0:4096-1];

  always @(posedge CLK) begin
    if(ram_w8_l16384_id2_0_0_enable) begin
      if(ram_w8_l16384_id2_0_0_wenable) begin
        mem[ram_w8_l16384_id2_0_0_addr] <= ram_w8_l16384_id2_0_0_wdata;
        ram_w8_l16384_id2_0_0_rdata_out <= ram_w8_l16384_id2_0_0_wdata;
      end else begin
        ram_w8_l16384_id2_0_0_rdata_out <= mem[ram_w8_l16384_id2_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l16384_id2_0_1_enable) begin
      if(ram_w8_l16384_id2_0_1_wenable) begin
        mem[ram_w8_l16384_id2_0_1_addr] <= ram_w8_l16384_id2_0_1_wdata;
        ram_w8_l16384_id2_0_1_rdata_out <= ram_w8_l16384_id2_0_1_wdata;
      end else begin
        ram_w8_l16384_id2_0_1_rdata_out <= mem[ram_w8_l16384_id2_0_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l16384_id2_1
(
  input CLK,
  input [12-1:0] ram_w8_l16384_id2_1_0_addr,
  output [8-1:0] ram_w8_l16384_id2_1_0_rdata,
  input [8-1:0] ram_w8_l16384_id2_1_0_wdata,
  input ram_w8_l16384_id2_1_0_wenable,
  input ram_w8_l16384_id2_1_0_enable,
  input [12-1:0] ram_w8_l16384_id2_1_1_addr,
  output [8-1:0] ram_w8_l16384_id2_1_1_rdata,
  input [8-1:0] ram_w8_l16384_id2_1_1_wdata,
  input ram_w8_l16384_id2_1_1_wenable,
  input ram_w8_l16384_id2_1_1_enable
);

  reg [8-1:0] ram_w8_l16384_id2_1_0_rdata_out;
  assign ram_w8_l16384_id2_1_0_rdata = ram_w8_l16384_id2_1_0_rdata_out;
  reg [8-1:0] ram_w8_l16384_id2_1_1_rdata_out;
  assign ram_w8_l16384_id2_1_1_rdata = ram_w8_l16384_id2_1_1_rdata_out;
  reg [8-1:0] mem [0:4096-1];

  always @(posedge CLK) begin
    if(ram_w8_l16384_id2_1_0_enable) begin
      if(ram_w8_l16384_id2_1_0_wenable) begin
        mem[ram_w8_l16384_id2_1_0_addr] <= ram_w8_l16384_id2_1_0_wdata;
        ram_w8_l16384_id2_1_0_rdata_out <= ram_w8_l16384_id2_1_0_wdata;
      end else begin
        ram_w8_l16384_id2_1_0_rdata_out <= mem[ram_w8_l16384_id2_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l16384_id2_1_1_enable) begin
      if(ram_w8_l16384_id2_1_1_wenable) begin
        mem[ram_w8_l16384_id2_1_1_addr] <= ram_w8_l16384_id2_1_1_wdata;
        ram_w8_l16384_id2_1_1_rdata_out <= ram_w8_l16384_id2_1_1_wdata;
      end else begin
        ram_w8_l16384_id2_1_1_rdata_out <= mem[ram_w8_l16384_id2_1_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l16384_id2_2
(
  input CLK,
  input [12-1:0] ram_w8_l16384_id2_2_0_addr,
  output [8-1:0] ram_w8_l16384_id2_2_0_rdata,
  input [8-1:0] ram_w8_l16384_id2_2_0_wdata,
  input ram_w8_l16384_id2_2_0_wenable,
  input ram_w8_l16384_id2_2_0_enable,
  input [12-1:0] ram_w8_l16384_id2_2_1_addr,
  output [8-1:0] ram_w8_l16384_id2_2_1_rdata,
  input [8-1:0] ram_w8_l16384_id2_2_1_wdata,
  input ram_w8_l16384_id2_2_1_wenable,
  input ram_w8_l16384_id2_2_1_enable
);

  reg [8-1:0] ram_w8_l16384_id2_2_0_rdata_out;
  assign ram_w8_l16384_id2_2_0_rdata = ram_w8_l16384_id2_2_0_rdata_out;
  reg [8-1:0] ram_w8_l16384_id2_2_1_rdata_out;
  assign ram_w8_l16384_id2_2_1_rdata = ram_w8_l16384_id2_2_1_rdata_out;
  reg [8-1:0] mem [0:4096-1];

  always @(posedge CLK) begin
    if(ram_w8_l16384_id2_2_0_enable) begin
      if(ram_w8_l16384_id2_2_0_wenable) begin
        mem[ram_w8_l16384_id2_2_0_addr] <= ram_w8_l16384_id2_2_0_wdata;
        ram_w8_l16384_id2_2_0_rdata_out <= ram_w8_l16384_id2_2_0_wdata;
      end else begin
        ram_w8_l16384_id2_2_0_rdata_out <= mem[ram_w8_l16384_id2_2_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l16384_id2_2_1_enable) begin
      if(ram_w8_l16384_id2_2_1_wenable) begin
        mem[ram_w8_l16384_id2_2_1_addr] <= ram_w8_l16384_id2_2_1_wdata;
        ram_w8_l16384_id2_2_1_rdata_out <= ram_w8_l16384_id2_2_1_wdata;
      end else begin
        ram_w8_l16384_id2_2_1_rdata_out <= mem[ram_w8_l16384_id2_2_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l16384_id2_3
(
  input CLK,
  input [12-1:0] ram_w8_l16384_id2_3_0_addr,
  output [8-1:0] ram_w8_l16384_id2_3_0_rdata,
  input [8-1:0] ram_w8_l16384_id2_3_0_wdata,
  input ram_w8_l16384_id2_3_0_wenable,
  input ram_w8_l16384_id2_3_0_enable,
  input [12-1:0] ram_w8_l16384_id2_3_1_addr,
  output [8-1:0] ram_w8_l16384_id2_3_1_rdata,
  input [8-1:0] ram_w8_l16384_id2_3_1_wdata,
  input ram_w8_l16384_id2_3_1_wenable,
  input ram_w8_l16384_id2_3_1_enable
);

  reg [8-1:0] ram_w8_l16384_id2_3_0_rdata_out;
  assign ram_w8_l16384_id2_3_0_rdata = ram_w8_l16384_id2_3_0_rdata_out;
  reg [8-1:0] ram_w8_l16384_id2_3_1_rdata_out;
  assign ram_w8_l16384_id2_3_1_rdata = ram_w8_l16384_id2_3_1_rdata_out;
  reg [8-1:0] mem [0:4096-1];

  always @(posedge CLK) begin
    if(ram_w8_l16384_id2_3_0_enable) begin
      if(ram_w8_l16384_id2_3_0_wenable) begin
        mem[ram_w8_l16384_id2_3_0_addr] <= ram_w8_l16384_id2_3_0_wdata;
        ram_w8_l16384_id2_3_0_rdata_out <= ram_w8_l16384_id2_3_0_wdata;
      end else begin
        ram_w8_l16384_id2_3_0_rdata_out <= mem[ram_w8_l16384_id2_3_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l16384_id2_3_1_enable) begin
      if(ram_w8_l16384_id2_3_1_wenable) begin
        mem[ram_w8_l16384_id2_3_1_addr] <= ram_w8_l16384_id2_3_1_wdata;
        ram_w8_l16384_id2_3_1_rdata_out <= ram_w8_l16384_id2_3_1_wdata;
      end else begin
        ram_w8_l16384_id2_3_1_rdata_out <= mem[ram_w8_l16384_id2_3_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l16384_id3_0
(
  input CLK,
  input [12-1:0] ram_w8_l16384_id3_0_0_addr,
  output [8-1:0] ram_w8_l16384_id3_0_0_rdata,
  input [8-1:0] ram_w8_l16384_id3_0_0_wdata,
  input ram_w8_l16384_id3_0_0_wenable,
  input ram_w8_l16384_id3_0_0_enable,
  input [12-1:0] ram_w8_l16384_id3_0_1_addr,
  output [8-1:0] ram_w8_l16384_id3_0_1_rdata,
  input [8-1:0] ram_w8_l16384_id3_0_1_wdata,
  input ram_w8_l16384_id3_0_1_wenable,
  input ram_w8_l16384_id3_0_1_enable
);

  reg [8-1:0] ram_w8_l16384_id3_0_0_rdata_out;
  assign ram_w8_l16384_id3_0_0_rdata = ram_w8_l16384_id3_0_0_rdata_out;
  reg [8-1:0] ram_w8_l16384_id3_0_1_rdata_out;
  assign ram_w8_l16384_id3_0_1_rdata = ram_w8_l16384_id3_0_1_rdata_out;
  reg [8-1:0] mem [0:4096-1];

  always @(posedge CLK) begin
    if(ram_w8_l16384_id3_0_0_enable) begin
      if(ram_w8_l16384_id3_0_0_wenable) begin
        mem[ram_w8_l16384_id3_0_0_addr] <= ram_w8_l16384_id3_0_0_wdata;
        ram_w8_l16384_id3_0_0_rdata_out <= ram_w8_l16384_id3_0_0_wdata;
      end else begin
        ram_w8_l16384_id3_0_0_rdata_out <= mem[ram_w8_l16384_id3_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l16384_id3_0_1_enable) begin
      if(ram_w8_l16384_id3_0_1_wenable) begin
        mem[ram_w8_l16384_id3_0_1_addr] <= ram_w8_l16384_id3_0_1_wdata;
        ram_w8_l16384_id3_0_1_rdata_out <= ram_w8_l16384_id3_0_1_wdata;
      end else begin
        ram_w8_l16384_id3_0_1_rdata_out <= mem[ram_w8_l16384_id3_0_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l16384_id3_1
(
  input CLK,
  input [12-1:0] ram_w8_l16384_id3_1_0_addr,
  output [8-1:0] ram_w8_l16384_id3_1_0_rdata,
  input [8-1:0] ram_w8_l16384_id3_1_0_wdata,
  input ram_w8_l16384_id3_1_0_wenable,
  input ram_w8_l16384_id3_1_0_enable,
  input [12-1:0] ram_w8_l16384_id3_1_1_addr,
  output [8-1:0] ram_w8_l16384_id3_1_1_rdata,
  input [8-1:0] ram_w8_l16384_id3_1_1_wdata,
  input ram_w8_l16384_id3_1_1_wenable,
  input ram_w8_l16384_id3_1_1_enable
);

  reg [8-1:0] ram_w8_l16384_id3_1_0_rdata_out;
  assign ram_w8_l16384_id3_1_0_rdata = ram_w8_l16384_id3_1_0_rdata_out;
  reg [8-1:0] ram_w8_l16384_id3_1_1_rdata_out;
  assign ram_w8_l16384_id3_1_1_rdata = ram_w8_l16384_id3_1_1_rdata_out;
  reg [8-1:0] mem [0:4096-1];

  always @(posedge CLK) begin
    if(ram_w8_l16384_id3_1_0_enable) begin
      if(ram_w8_l16384_id3_1_0_wenable) begin
        mem[ram_w8_l16384_id3_1_0_addr] <= ram_w8_l16384_id3_1_0_wdata;
        ram_w8_l16384_id3_1_0_rdata_out <= ram_w8_l16384_id3_1_0_wdata;
      end else begin
        ram_w8_l16384_id3_1_0_rdata_out <= mem[ram_w8_l16384_id3_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l16384_id3_1_1_enable) begin
      if(ram_w8_l16384_id3_1_1_wenable) begin
        mem[ram_w8_l16384_id3_1_1_addr] <= ram_w8_l16384_id3_1_1_wdata;
        ram_w8_l16384_id3_1_1_rdata_out <= ram_w8_l16384_id3_1_1_wdata;
      end else begin
        ram_w8_l16384_id3_1_1_rdata_out <= mem[ram_w8_l16384_id3_1_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l16384_id3_2
(
  input CLK,
  input [12-1:0] ram_w8_l16384_id3_2_0_addr,
  output [8-1:0] ram_w8_l16384_id3_2_0_rdata,
  input [8-1:0] ram_w8_l16384_id3_2_0_wdata,
  input ram_w8_l16384_id3_2_0_wenable,
  input ram_w8_l16384_id3_2_0_enable,
  input [12-1:0] ram_w8_l16384_id3_2_1_addr,
  output [8-1:0] ram_w8_l16384_id3_2_1_rdata,
  input [8-1:0] ram_w8_l16384_id3_2_1_wdata,
  input ram_w8_l16384_id3_2_1_wenable,
  input ram_w8_l16384_id3_2_1_enable
);

  reg [8-1:0] ram_w8_l16384_id3_2_0_rdata_out;
  assign ram_w8_l16384_id3_2_0_rdata = ram_w8_l16384_id3_2_0_rdata_out;
  reg [8-1:0] ram_w8_l16384_id3_2_1_rdata_out;
  assign ram_w8_l16384_id3_2_1_rdata = ram_w8_l16384_id3_2_1_rdata_out;
  reg [8-1:0] mem [0:4096-1];

  always @(posedge CLK) begin
    if(ram_w8_l16384_id3_2_0_enable) begin
      if(ram_w8_l16384_id3_2_0_wenable) begin
        mem[ram_w8_l16384_id3_2_0_addr] <= ram_w8_l16384_id3_2_0_wdata;
        ram_w8_l16384_id3_2_0_rdata_out <= ram_w8_l16384_id3_2_0_wdata;
      end else begin
        ram_w8_l16384_id3_2_0_rdata_out <= mem[ram_w8_l16384_id3_2_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l16384_id3_2_1_enable) begin
      if(ram_w8_l16384_id3_2_1_wenable) begin
        mem[ram_w8_l16384_id3_2_1_addr] <= ram_w8_l16384_id3_2_1_wdata;
        ram_w8_l16384_id3_2_1_rdata_out <= ram_w8_l16384_id3_2_1_wdata;
      end else begin
        ram_w8_l16384_id3_2_1_rdata_out <= mem[ram_w8_l16384_id3_2_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l16384_id3_3
(
  input CLK,
  input [12-1:0] ram_w8_l16384_id3_3_0_addr,
  output [8-1:0] ram_w8_l16384_id3_3_0_rdata,
  input [8-1:0] ram_w8_l16384_id3_3_0_wdata,
  input ram_w8_l16384_id3_3_0_wenable,
  input ram_w8_l16384_id3_3_0_enable,
  input [12-1:0] ram_w8_l16384_id3_3_1_addr,
  output [8-1:0] ram_w8_l16384_id3_3_1_rdata,
  input [8-1:0] ram_w8_l16384_id3_3_1_wdata,
  input ram_w8_l16384_id3_3_1_wenable,
  input ram_w8_l16384_id3_3_1_enable
);

  reg [8-1:0] ram_w8_l16384_id3_3_0_rdata_out;
  assign ram_w8_l16384_id3_3_0_rdata = ram_w8_l16384_id3_3_0_rdata_out;
  reg [8-1:0] ram_w8_l16384_id3_3_1_rdata_out;
  assign ram_w8_l16384_id3_3_1_rdata = ram_w8_l16384_id3_3_1_rdata_out;
  reg [8-1:0] mem [0:4096-1];

  always @(posedge CLK) begin
    if(ram_w8_l16384_id3_3_0_enable) begin
      if(ram_w8_l16384_id3_3_0_wenable) begin
        mem[ram_w8_l16384_id3_3_0_addr] <= ram_w8_l16384_id3_3_0_wdata;
        ram_w8_l16384_id3_3_0_rdata_out <= ram_w8_l16384_id3_3_0_wdata;
      end else begin
        ram_w8_l16384_id3_3_0_rdata_out <= mem[ram_w8_l16384_id3_3_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l16384_id3_3_1_enable) begin
      if(ram_w8_l16384_id3_3_1_wenable) begin
        mem[ram_w8_l16384_id3_3_1_addr] <= ram_w8_l16384_id3_3_1_wdata;
        ram_w8_l16384_id3_3_1_rdata_out <= ram_w8_l16384_id3_3_1_wdata;
      end else begin
        ram_w8_l16384_id3_3_1_rdata_out <= mem[ram_w8_l16384_id3_3_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l16384_id4_0
(
  input CLK,
  input [12-1:0] ram_w8_l16384_id4_0_0_addr,
  output [8-1:0] ram_w8_l16384_id4_0_0_rdata,
  input [8-1:0] ram_w8_l16384_id4_0_0_wdata,
  input ram_w8_l16384_id4_0_0_wenable,
  input ram_w8_l16384_id4_0_0_enable,
  input [12-1:0] ram_w8_l16384_id4_0_1_addr,
  output [8-1:0] ram_w8_l16384_id4_0_1_rdata,
  input [8-1:0] ram_w8_l16384_id4_0_1_wdata,
  input ram_w8_l16384_id4_0_1_wenable,
  input ram_w8_l16384_id4_0_1_enable
);

  reg [8-1:0] ram_w8_l16384_id4_0_0_rdata_out;
  assign ram_w8_l16384_id4_0_0_rdata = ram_w8_l16384_id4_0_0_rdata_out;
  reg [8-1:0] ram_w8_l16384_id4_0_1_rdata_out;
  assign ram_w8_l16384_id4_0_1_rdata = ram_w8_l16384_id4_0_1_rdata_out;
  reg [8-1:0] mem [0:4096-1];

  always @(posedge CLK) begin
    if(ram_w8_l16384_id4_0_0_enable) begin
      if(ram_w8_l16384_id4_0_0_wenable) begin
        mem[ram_w8_l16384_id4_0_0_addr] <= ram_w8_l16384_id4_0_0_wdata;
        ram_w8_l16384_id4_0_0_rdata_out <= ram_w8_l16384_id4_0_0_wdata;
      end else begin
        ram_w8_l16384_id4_0_0_rdata_out <= mem[ram_w8_l16384_id4_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l16384_id4_0_1_enable) begin
      if(ram_w8_l16384_id4_0_1_wenable) begin
        mem[ram_w8_l16384_id4_0_1_addr] <= ram_w8_l16384_id4_0_1_wdata;
        ram_w8_l16384_id4_0_1_rdata_out <= ram_w8_l16384_id4_0_1_wdata;
      end else begin
        ram_w8_l16384_id4_0_1_rdata_out <= mem[ram_w8_l16384_id4_0_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l16384_id4_1
(
  input CLK,
  input [12-1:0] ram_w8_l16384_id4_1_0_addr,
  output [8-1:0] ram_w8_l16384_id4_1_0_rdata,
  input [8-1:0] ram_w8_l16384_id4_1_0_wdata,
  input ram_w8_l16384_id4_1_0_wenable,
  input ram_w8_l16384_id4_1_0_enable,
  input [12-1:0] ram_w8_l16384_id4_1_1_addr,
  output [8-1:0] ram_w8_l16384_id4_1_1_rdata,
  input [8-1:0] ram_w8_l16384_id4_1_1_wdata,
  input ram_w8_l16384_id4_1_1_wenable,
  input ram_w8_l16384_id4_1_1_enable
);

  reg [8-1:0] ram_w8_l16384_id4_1_0_rdata_out;
  assign ram_w8_l16384_id4_1_0_rdata = ram_w8_l16384_id4_1_0_rdata_out;
  reg [8-1:0] ram_w8_l16384_id4_1_1_rdata_out;
  assign ram_w8_l16384_id4_1_1_rdata = ram_w8_l16384_id4_1_1_rdata_out;
  reg [8-1:0] mem [0:4096-1];

  always @(posedge CLK) begin
    if(ram_w8_l16384_id4_1_0_enable) begin
      if(ram_w8_l16384_id4_1_0_wenable) begin
        mem[ram_w8_l16384_id4_1_0_addr] <= ram_w8_l16384_id4_1_0_wdata;
        ram_w8_l16384_id4_1_0_rdata_out <= ram_w8_l16384_id4_1_0_wdata;
      end else begin
        ram_w8_l16384_id4_1_0_rdata_out <= mem[ram_w8_l16384_id4_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l16384_id4_1_1_enable) begin
      if(ram_w8_l16384_id4_1_1_wenable) begin
        mem[ram_w8_l16384_id4_1_1_addr] <= ram_w8_l16384_id4_1_1_wdata;
        ram_w8_l16384_id4_1_1_rdata_out <= ram_w8_l16384_id4_1_1_wdata;
      end else begin
        ram_w8_l16384_id4_1_1_rdata_out <= mem[ram_w8_l16384_id4_1_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l16384_id4_2
(
  input CLK,
  input [12-1:0] ram_w8_l16384_id4_2_0_addr,
  output [8-1:0] ram_w8_l16384_id4_2_0_rdata,
  input [8-1:0] ram_w8_l16384_id4_2_0_wdata,
  input ram_w8_l16384_id4_2_0_wenable,
  input ram_w8_l16384_id4_2_0_enable,
  input [12-1:0] ram_w8_l16384_id4_2_1_addr,
  output [8-1:0] ram_w8_l16384_id4_2_1_rdata,
  input [8-1:0] ram_w8_l16384_id4_2_1_wdata,
  input ram_w8_l16384_id4_2_1_wenable,
  input ram_w8_l16384_id4_2_1_enable
);

  reg [8-1:0] ram_w8_l16384_id4_2_0_rdata_out;
  assign ram_w8_l16384_id4_2_0_rdata = ram_w8_l16384_id4_2_0_rdata_out;
  reg [8-1:0] ram_w8_l16384_id4_2_1_rdata_out;
  assign ram_w8_l16384_id4_2_1_rdata = ram_w8_l16384_id4_2_1_rdata_out;
  reg [8-1:0] mem [0:4096-1];

  always @(posedge CLK) begin
    if(ram_w8_l16384_id4_2_0_enable) begin
      if(ram_w8_l16384_id4_2_0_wenable) begin
        mem[ram_w8_l16384_id4_2_0_addr] <= ram_w8_l16384_id4_2_0_wdata;
        ram_w8_l16384_id4_2_0_rdata_out <= ram_w8_l16384_id4_2_0_wdata;
      end else begin
        ram_w8_l16384_id4_2_0_rdata_out <= mem[ram_w8_l16384_id4_2_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l16384_id4_2_1_enable) begin
      if(ram_w8_l16384_id4_2_1_wenable) begin
        mem[ram_w8_l16384_id4_2_1_addr] <= ram_w8_l16384_id4_2_1_wdata;
        ram_w8_l16384_id4_2_1_rdata_out <= ram_w8_l16384_id4_2_1_wdata;
      end else begin
        ram_w8_l16384_id4_2_1_rdata_out <= mem[ram_w8_l16384_id4_2_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l16384_id4_3
(
  input CLK,
  input [12-1:0] ram_w8_l16384_id4_3_0_addr,
  output [8-1:0] ram_w8_l16384_id4_3_0_rdata,
  input [8-1:0] ram_w8_l16384_id4_3_0_wdata,
  input ram_w8_l16384_id4_3_0_wenable,
  input ram_w8_l16384_id4_3_0_enable,
  input [12-1:0] ram_w8_l16384_id4_3_1_addr,
  output [8-1:0] ram_w8_l16384_id4_3_1_rdata,
  input [8-1:0] ram_w8_l16384_id4_3_1_wdata,
  input ram_w8_l16384_id4_3_1_wenable,
  input ram_w8_l16384_id4_3_1_enable
);

  reg [8-1:0] ram_w8_l16384_id4_3_0_rdata_out;
  assign ram_w8_l16384_id4_3_0_rdata = ram_w8_l16384_id4_3_0_rdata_out;
  reg [8-1:0] ram_w8_l16384_id4_3_1_rdata_out;
  assign ram_w8_l16384_id4_3_1_rdata = ram_w8_l16384_id4_3_1_rdata_out;
  reg [8-1:0] mem [0:4096-1];

  always @(posedge CLK) begin
    if(ram_w8_l16384_id4_3_0_enable) begin
      if(ram_w8_l16384_id4_3_0_wenable) begin
        mem[ram_w8_l16384_id4_3_0_addr] <= ram_w8_l16384_id4_3_0_wdata;
        ram_w8_l16384_id4_3_0_rdata_out <= ram_w8_l16384_id4_3_0_wdata;
      end else begin
        ram_w8_l16384_id4_3_0_rdata_out <= mem[ram_w8_l16384_id4_3_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l16384_id4_3_1_enable) begin
      if(ram_w8_l16384_id4_3_1_wenable) begin
        mem[ram_w8_l16384_id4_3_1_addr] <= ram_w8_l16384_id4_3_1_wdata;
        ram_w8_l16384_id4_3_1_rdata_out <= ram_w8_l16384_id4_3_1_wdata;
      end else begin
        ram_w8_l16384_id4_3_1_rdata_out <= mem[ram_w8_l16384_id4_3_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l16384_id5_0
(
  input CLK,
  input [12-1:0] ram_w8_l16384_id5_0_0_addr,
  output [8-1:0] ram_w8_l16384_id5_0_0_rdata,
  input [8-1:0] ram_w8_l16384_id5_0_0_wdata,
  input ram_w8_l16384_id5_0_0_wenable,
  input ram_w8_l16384_id5_0_0_enable,
  input [12-1:0] ram_w8_l16384_id5_0_1_addr,
  output [8-1:0] ram_w8_l16384_id5_0_1_rdata,
  input [8-1:0] ram_w8_l16384_id5_0_1_wdata,
  input ram_w8_l16384_id5_0_1_wenable,
  input ram_w8_l16384_id5_0_1_enable
);

  reg [8-1:0] ram_w8_l16384_id5_0_0_rdata_out;
  assign ram_w8_l16384_id5_0_0_rdata = ram_w8_l16384_id5_0_0_rdata_out;
  reg [8-1:0] ram_w8_l16384_id5_0_1_rdata_out;
  assign ram_w8_l16384_id5_0_1_rdata = ram_w8_l16384_id5_0_1_rdata_out;
  reg [8-1:0] mem [0:4096-1];

  always @(posedge CLK) begin
    if(ram_w8_l16384_id5_0_0_enable) begin
      if(ram_w8_l16384_id5_0_0_wenable) begin
        mem[ram_w8_l16384_id5_0_0_addr] <= ram_w8_l16384_id5_0_0_wdata;
        ram_w8_l16384_id5_0_0_rdata_out <= ram_w8_l16384_id5_0_0_wdata;
      end else begin
        ram_w8_l16384_id5_0_0_rdata_out <= mem[ram_w8_l16384_id5_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l16384_id5_0_1_enable) begin
      if(ram_w8_l16384_id5_0_1_wenable) begin
        mem[ram_w8_l16384_id5_0_1_addr] <= ram_w8_l16384_id5_0_1_wdata;
        ram_w8_l16384_id5_0_1_rdata_out <= ram_w8_l16384_id5_0_1_wdata;
      end else begin
        ram_w8_l16384_id5_0_1_rdata_out <= mem[ram_w8_l16384_id5_0_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l16384_id5_1
(
  input CLK,
  input [12-1:0] ram_w8_l16384_id5_1_0_addr,
  output [8-1:0] ram_w8_l16384_id5_1_0_rdata,
  input [8-1:0] ram_w8_l16384_id5_1_0_wdata,
  input ram_w8_l16384_id5_1_0_wenable,
  input ram_w8_l16384_id5_1_0_enable,
  input [12-1:0] ram_w8_l16384_id5_1_1_addr,
  output [8-1:0] ram_w8_l16384_id5_1_1_rdata,
  input [8-1:0] ram_w8_l16384_id5_1_1_wdata,
  input ram_w8_l16384_id5_1_1_wenable,
  input ram_w8_l16384_id5_1_1_enable
);

  reg [8-1:0] ram_w8_l16384_id5_1_0_rdata_out;
  assign ram_w8_l16384_id5_1_0_rdata = ram_w8_l16384_id5_1_0_rdata_out;
  reg [8-1:0] ram_w8_l16384_id5_1_1_rdata_out;
  assign ram_w8_l16384_id5_1_1_rdata = ram_w8_l16384_id5_1_1_rdata_out;
  reg [8-1:0] mem [0:4096-1];

  always @(posedge CLK) begin
    if(ram_w8_l16384_id5_1_0_enable) begin
      if(ram_w8_l16384_id5_1_0_wenable) begin
        mem[ram_w8_l16384_id5_1_0_addr] <= ram_w8_l16384_id5_1_0_wdata;
        ram_w8_l16384_id5_1_0_rdata_out <= ram_w8_l16384_id5_1_0_wdata;
      end else begin
        ram_w8_l16384_id5_1_0_rdata_out <= mem[ram_w8_l16384_id5_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l16384_id5_1_1_enable) begin
      if(ram_w8_l16384_id5_1_1_wenable) begin
        mem[ram_w8_l16384_id5_1_1_addr] <= ram_w8_l16384_id5_1_1_wdata;
        ram_w8_l16384_id5_1_1_rdata_out <= ram_w8_l16384_id5_1_1_wdata;
      end else begin
        ram_w8_l16384_id5_1_1_rdata_out <= mem[ram_w8_l16384_id5_1_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l16384_id5_2
(
  input CLK,
  input [12-1:0] ram_w8_l16384_id5_2_0_addr,
  output [8-1:0] ram_w8_l16384_id5_2_0_rdata,
  input [8-1:0] ram_w8_l16384_id5_2_0_wdata,
  input ram_w8_l16384_id5_2_0_wenable,
  input ram_w8_l16384_id5_2_0_enable,
  input [12-1:0] ram_w8_l16384_id5_2_1_addr,
  output [8-1:0] ram_w8_l16384_id5_2_1_rdata,
  input [8-1:0] ram_w8_l16384_id5_2_1_wdata,
  input ram_w8_l16384_id5_2_1_wenable,
  input ram_w8_l16384_id5_2_1_enable
);

  reg [8-1:0] ram_w8_l16384_id5_2_0_rdata_out;
  assign ram_w8_l16384_id5_2_0_rdata = ram_w8_l16384_id5_2_0_rdata_out;
  reg [8-1:0] ram_w8_l16384_id5_2_1_rdata_out;
  assign ram_w8_l16384_id5_2_1_rdata = ram_w8_l16384_id5_2_1_rdata_out;
  reg [8-1:0] mem [0:4096-1];

  always @(posedge CLK) begin
    if(ram_w8_l16384_id5_2_0_enable) begin
      if(ram_w8_l16384_id5_2_0_wenable) begin
        mem[ram_w8_l16384_id5_2_0_addr] <= ram_w8_l16384_id5_2_0_wdata;
        ram_w8_l16384_id5_2_0_rdata_out <= ram_w8_l16384_id5_2_0_wdata;
      end else begin
        ram_w8_l16384_id5_2_0_rdata_out <= mem[ram_w8_l16384_id5_2_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l16384_id5_2_1_enable) begin
      if(ram_w8_l16384_id5_2_1_wenable) begin
        mem[ram_w8_l16384_id5_2_1_addr] <= ram_w8_l16384_id5_2_1_wdata;
        ram_w8_l16384_id5_2_1_rdata_out <= ram_w8_l16384_id5_2_1_wdata;
      end else begin
        ram_w8_l16384_id5_2_1_rdata_out <= mem[ram_w8_l16384_id5_2_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l16384_id5_3
(
  input CLK,
  input [12-1:0] ram_w8_l16384_id5_3_0_addr,
  output [8-1:0] ram_w8_l16384_id5_3_0_rdata,
  input [8-1:0] ram_w8_l16384_id5_3_0_wdata,
  input ram_w8_l16384_id5_3_0_wenable,
  input ram_w8_l16384_id5_3_0_enable,
  input [12-1:0] ram_w8_l16384_id5_3_1_addr,
  output [8-1:0] ram_w8_l16384_id5_3_1_rdata,
  input [8-1:0] ram_w8_l16384_id5_3_1_wdata,
  input ram_w8_l16384_id5_3_1_wenable,
  input ram_w8_l16384_id5_3_1_enable
);

  reg [8-1:0] ram_w8_l16384_id5_3_0_rdata_out;
  assign ram_w8_l16384_id5_3_0_rdata = ram_w8_l16384_id5_3_0_rdata_out;
  reg [8-1:0] ram_w8_l16384_id5_3_1_rdata_out;
  assign ram_w8_l16384_id5_3_1_rdata = ram_w8_l16384_id5_3_1_rdata_out;
  reg [8-1:0] mem [0:4096-1];

  always @(posedge CLK) begin
    if(ram_w8_l16384_id5_3_0_enable) begin
      if(ram_w8_l16384_id5_3_0_wenable) begin
        mem[ram_w8_l16384_id5_3_0_addr] <= ram_w8_l16384_id5_3_0_wdata;
        ram_w8_l16384_id5_3_0_rdata_out <= ram_w8_l16384_id5_3_0_wdata;
      end else begin
        ram_w8_l16384_id5_3_0_rdata_out <= mem[ram_w8_l16384_id5_3_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l16384_id5_3_1_enable) begin
      if(ram_w8_l16384_id5_3_1_wenable) begin
        mem[ram_w8_l16384_id5_3_1_addr] <= ram_w8_l16384_id5_3_1_wdata;
        ram_w8_l16384_id5_3_1_rdata_out <= ram_w8_l16384_id5_3_1_wdata;
      end else begin
        ram_w8_l16384_id5_3_1_rdata_out <= mem[ram_w8_l16384_id5_3_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l16384_id6_0
(
  input CLK,
  input [12-1:0] ram_w8_l16384_id6_0_0_addr,
  output [8-1:0] ram_w8_l16384_id6_0_0_rdata,
  input [8-1:0] ram_w8_l16384_id6_0_0_wdata,
  input ram_w8_l16384_id6_0_0_wenable,
  input ram_w8_l16384_id6_0_0_enable,
  input [12-1:0] ram_w8_l16384_id6_0_1_addr,
  output [8-1:0] ram_w8_l16384_id6_0_1_rdata,
  input [8-1:0] ram_w8_l16384_id6_0_1_wdata,
  input ram_w8_l16384_id6_0_1_wenable,
  input ram_w8_l16384_id6_0_1_enable
);

  reg [8-1:0] ram_w8_l16384_id6_0_0_rdata_out;
  assign ram_w8_l16384_id6_0_0_rdata = ram_w8_l16384_id6_0_0_rdata_out;
  reg [8-1:0] ram_w8_l16384_id6_0_1_rdata_out;
  assign ram_w8_l16384_id6_0_1_rdata = ram_w8_l16384_id6_0_1_rdata_out;
  reg [8-1:0] mem [0:4096-1];

  always @(posedge CLK) begin
    if(ram_w8_l16384_id6_0_0_enable) begin
      if(ram_w8_l16384_id6_0_0_wenable) begin
        mem[ram_w8_l16384_id6_0_0_addr] <= ram_w8_l16384_id6_0_0_wdata;
        ram_w8_l16384_id6_0_0_rdata_out <= ram_w8_l16384_id6_0_0_wdata;
      end else begin
        ram_w8_l16384_id6_0_0_rdata_out <= mem[ram_w8_l16384_id6_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l16384_id6_0_1_enable) begin
      if(ram_w8_l16384_id6_0_1_wenable) begin
        mem[ram_w8_l16384_id6_0_1_addr] <= ram_w8_l16384_id6_0_1_wdata;
        ram_w8_l16384_id6_0_1_rdata_out <= ram_w8_l16384_id6_0_1_wdata;
      end else begin
        ram_w8_l16384_id6_0_1_rdata_out <= mem[ram_w8_l16384_id6_0_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l16384_id6_1
(
  input CLK,
  input [12-1:0] ram_w8_l16384_id6_1_0_addr,
  output [8-1:0] ram_w8_l16384_id6_1_0_rdata,
  input [8-1:0] ram_w8_l16384_id6_1_0_wdata,
  input ram_w8_l16384_id6_1_0_wenable,
  input ram_w8_l16384_id6_1_0_enable,
  input [12-1:0] ram_w8_l16384_id6_1_1_addr,
  output [8-1:0] ram_w8_l16384_id6_1_1_rdata,
  input [8-1:0] ram_w8_l16384_id6_1_1_wdata,
  input ram_w8_l16384_id6_1_1_wenable,
  input ram_w8_l16384_id6_1_1_enable
);

  reg [8-1:0] ram_w8_l16384_id6_1_0_rdata_out;
  assign ram_w8_l16384_id6_1_0_rdata = ram_w8_l16384_id6_1_0_rdata_out;
  reg [8-1:0] ram_w8_l16384_id6_1_1_rdata_out;
  assign ram_w8_l16384_id6_1_1_rdata = ram_w8_l16384_id6_1_1_rdata_out;
  reg [8-1:0] mem [0:4096-1];

  always @(posedge CLK) begin
    if(ram_w8_l16384_id6_1_0_enable) begin
      if(ram_w8_l16384_id6_1_0_wenable) begin
        mem[ram_w8_l16384_id6_1_0_addr] <= ram_w8_l16384_id6_1_0_wdata;
        ram_w8_l16384_id6_1_0_rdata_out <= ram_w8_l16384_id6_1_0_wdata;
      end else begin
        ram_w8_l16384_id6_1_0_rdata_out <= mem[ram_w8_l16384_id6_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l16384_id6_1_1_enable) begin
      if(ram_w8_l16384_id6_1_1_wenable) begin
        mem[ram_w8_l16384_id6_1_1_addr] <= ram_w8_l16384_id6_1_1_wdata;
        ram_w8_l16384_id6_1_1_rdata_out <= ram_w8_l16384_id6_1_1_wdata;
      end else begin
        ram_w8_l16384_id6_1_1_rdata_out <= mem[ram_w8_l16384_id6_1_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l16384_id6_2
(
  input CLK,
  input [12-1:0] ram_w8_l16384_id6_2_0_addr,
  output [8-1:0] ram_w8_l16384_id6_2_0_rdata,
  input [8-1:0] ram_w8_l16384_id6_2_0_wdata,
  input ram_w8_l16384_id6_2_0_wenable,
  input ram_w8_l16384_id6_2_0_enable,
  input [12-1:0] ram_w8_l16384_id6_2_1_addr,
  output [8-1:0] ram_w8_l16384_id6_2_1_rdata,
  input [8-1:0] ram_w8_l16384_id6_2_1_wdata,
  input ram_w8_l16384_id6_2_1_wenable,
  input ram_w8_l16384_id6_2_1_enable
);

  reg [8-1:0] ram_w8_l16384_id6_2_0_rdata_out;
  assign ram_w8_l16384_id6_2_0_rdata = ram_w8_l16384_id6_2_0_rdata_out;
  reg [8-1:0] ram_w8_l16384_id6_2_1_rdata_out;
  assign ram_w8_l16384_id6_2_1_rdata = ram_w8_l16384_id6_2_1_rdata_out;
  reg [8-1:0] mem [0:4096-1];

  always @(posedge CLK) begin
    if(ram_w8_l16384_id6_2_0_enable) begin
      if(ram_w8_l16384_id6_2_0_wenable) begin
        mem[ram_w8_l16384_id6_2_0_addr] <= ram_w8_l16384_id6_2_0_wdata;
        ram_w8_l16384_id6_2_0_rdata_out <= ram_w8_l16384_id6_2_0_wdata;
      end else begin
        ram_w8_l16384_id6_2_0_rdata_out <= mem[ram_w8_l16384_id6_2_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l16384_id6_2_1_enable) begin
      if(ram_w8_l16384_id6_2_1_wenable) begin
        mem[ram_w8_l16384_id6_2_1_addr] <= ram_w8_l16384_id6_2_1_wdata;
        ram_w8_l16384_id6_2_1_rdata_out <= ram_w8_l16384_id6_2_1_wdata;
      end else begin
        ram_w8_l16384_id6_2_1_rdata_out <= mem[ram_w8_l16384_id6_2_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l16384_id6_3
(
  input CLK,
  input [12-1:0] ram_w8_l16384_id6_3_0_addr,
  output [8-1:0] ram_w8_l16384_id6_3_0_rdata,
  input [8-1:0] ram_w8_l16384_id6_3_0_wdata,
  input ram_w8_l16384_id6_3_0_wenable,
  input ram_w8_l16384_id6_3_0_enable,
  input [12-1:0] ram_w8_l16384_id6_3_1_addr,
  output [8-1:0] ram_w8_l16384_id6_3_1_rdata,
  input [8-1:0] ram_w8_l16384_id6_3_1_wdata,
  input ram_w8_l16384_id6_3_1_wenable,
  input ram_w8_l16384_id6_3_1_enable
);

  reg [8-1:0] ram_w8_l16384_id6_3_0_rdata_out;
  assign ram_w8_l16384_id6_3_0_rdata = ram_w8_l16384_id6_3_0_rdata_out;
  reg [8-1:0] ram_w8_l16384_id6_3_1_rdata_out;
  assign ram_w8_l16384_id6_3_1_rdata = ram_w8_l16384_id6_3_1_rdata_out;
  reg [8-1:0] mem [0:4096-1];

  always @(posedge CLK) begin
    if(ram_w8_l16384_id6_3_0_enable) begin
      if(ram_w8_l16384_id6_3_0_wenable) begin
        mem[ram_w8_l16384_id6_3_0_addr] <= ram_w8_l16384_id6_3_0_wdata;
        ram_w8_l16384_id6_3_0_rdata_out <= ram_w8_l16384_id6_3_0_wdata;
      end else begin
        ram_w8_l16384_id6_3_0_rdata_out <= mem[ram_w8_l16384_id6_3_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l16384_id6_3_1_enable) begin
      if(ram_w8_l16384_id6_3_1_wenable) begin
        mem[ram_w8_l16384_id6_3_1_addr] <= ram_w8_l16384_id6_3_1_wdata;
        ram_w8_l16384_id6_3_1_rdata_out <= ram_w8_l16384_id6_3_1_wdata;
      end else begin
        ram_w8_l16384_id6_3_1_rdata_out <= mem[ram_w8_l16384_id6_3_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l16384_id7_0
(
  input CLK,
  input [12-1:0] ram_w8_l16384_id7_0_0_addr,
  output [8-1:0] ram_w8_l16384_id7_0_0_rdata,
  input [8-1:0] ram_w8_l16384_id7_0_0_wdata,
  input ram_w8_l16384_id7_0_0_wenable,
  input ram_w8_l16384_id7_0_0_enable,
  input [12-1:0] ram_w8_l16384_id7_0_1_addr,
  output [8-1:0] ram_w8_l16384_id7_0_1_rdata,
  input [8-1:0] ram_w8_l16384_id7_0_1_wdata,
  input ram_w8_l16384_id7_0_1_wenable,
  input ram_w8_l16384_id7_0_1_enable
);

  reg [8-1:0] ram_w8_l16384_id7_0_0_rdata_out;
  assign ram_w8_l16384_id7_0_0_rdata = ram_w8_l16384_id7_0_0_rdata_out;
  reg [8-1:0] ram_w8_l16384_id7_0_1_rdata_out;
  assign ram_w8_l16384_id7_0_1_rdata = ram_w8_l16384_id7_0_1_rdata_out;
  reg [8-1:0] mem [0:4096-1];

  always @(posedge CLK) begin
    if(ram_w8_l16384_id7_0_0_enable) begin
      if(ram_w8_l16384_id7_0_0_wenable) begin
        mem[ram_w8_l16384_id7_0_0_addr] <= ram_w8_l16384_id7_0_0_wdata;
        ram_w8_l16384_id7_0_0_rdata_out <= ram_w8_l16384_id7_0_0_wdata;
      end else begin
        ram_w8_l16384_id7_0_0_rdata_out <= mem[ram_w8_l16384_id7_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l16384_id7_0_1_enable) begin
      if(ram_w8_l16384_id7_0_1_wenable) begin
        mem[ram_w8_l16384_id7_0_1_addr] <= ram_w8_l16384_id7_0_1_wdata;
        ram_w8_l16384_id7_0_1_rdata_out <= ram_w8_l16384_id7_0_1_wdata;
      end else begin
        ram_w8_l16384_id7_0_1_rdata_out <= mem[ram_w8_l16384_id7_0_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l16384_id7_1
(
  input CLK,
  input [12-1:0] ram_w8_l16384_id7_1_0_addr,
  output [8-1:0] ram_w8_l16384_id7_1_0_rdata,
  input [8-1:0] ram_w8_l16384_id7_1_0_wdata,
  input ram_w8_l16384_id7_1_0_wenable,
  input ram_w8_l16384_id7_1_0_enable,
  input [12-1:0] ram_w8_l16384_id7_1_1_addr,
  output [8-1:0] ram_w8_l16384_id7_1_1_rdata,
  input [8-1:0] ram_w8_l16384_id7_1_1_wdata,
  input ram_w8_l16384_id7_1_1_wenable,
  input ram_w8_l16384_id7_1_1_enable
);

  reg [8-1:0] ram_w8_l16384_id7_1_0_rdata_out;
  assign ram_w8_l16384_id7_1_0_rdata = ram_w8_l16384_id7_1_0_rdata_out;
  reg [8-1:0] ram_w8_l16384_id7_1_1_rdata_out;
  assign ram_w8_l16384_id7_1_1_rdata = ram_w8_l16384_id7_1_1_rdata_out;
  reg [8-1:0] mem [0:4096-1];

  always @(posedge CLK) begin
    if(ram_w8_l16384_id7_1_0_enable) begin
      if(ram_w8_l16384_id7_1_0_wenable) begin
        mem[ram_w8_l16384_id7_1_0_addr] <= ram_w8_l16384_id7_1_0_wdata;
        ram_w8_l16384_id7_1_0_rdata_out <= ram_w8_l16384_id7_1_0_wdata;
      end else begin
        ram_w8_l16384_id7_1_0_rdata_out <= mem[ram_w8_l16384_id7_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l16384_id7_1_1_enable) begin
      if(ram_w8_l16384_id7_1_1_wenable) begin
        mem[ram_w8_l16384_id7_1_1_addr] <= ram_w8_l16384_id7_1_1_wdata;
        ram_w8_l16384_id7_1_1_rdata_out <= ram_w8_l16384_id7_1_1_wdata;
      end else begin
        ram_w8_l16384_id7_1_1_rdata_out <= mem[ram_w8_l16384_id7_1_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l16384_id7_2
(
  input CLK,
  input [12-1:0] ram_w8_l16384_id7_2_0_addr,
  output [8-1:0] ram_w8_l16384_id7_2_0_rdata,
  input [8-1:0] ram_w8_l16384_id7_2_0_wdata,
  input ram_w8_l16384_id7_2_0_wenable,
  input ram_w8_l16384_id7_2_0_enable,
  input [12-1:0] ram_w8_l16384_id7_2_1_addr,
  output [8-1:0] ram_w8_l16384_id7_2_1_rdata,
  input [8-1:0] ram_w8_l16384_id7_2_1_wdata,
  input ram_w8_l16384_id7_2_1_wenable,
  input ram_w8_l16384_id7_2_1_enable
);

  reg [8-1:0] ram_w8_l16384_id7_2_0_rdata_out;
  assign ram_w8_l16384_id7_2_0_rdata = ram_w8_l16384_id7_2_0_rdata_out;
  reg [8-1:0] ram_w8_l16384_id7_2_1_rdata_out;
  assign ram_w8_l16384_id7_2_1_rdata = ram_w8_l16384_id7_2_1_rdata_out;
  reg [8-1:0] mem [0:4096-1];

  always @(posedge CLK) begin
    if(ram_w8_l16384_id7_2_0_enable) begin
      if(ram_w8_l16384_id7_2_0_wenable) begin
        mem[ram_w8_l16384_id7_2_0_addr] <= ram_w8_l16384_id7_2_0_wdata;
        ram_w8_l16384_id7_2_0_rdata_out <= ram_w8_l16384_id7_2_0_wdata;
      end else begin
        ram_w8_l16384_id7_2_0_rdata_out <= mem[ram_w8_l16384_id7_2_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l16384_id7_2_1_enable) begin
      if(ram_w8_l16384_id7_2_1_wenable) begin
        mem[ram_w8_l16384_id7_2_1_addr] <= ram_w8_l16384_id7_2_1_wdata;
        ram_w8_l16384_id7_2_1_rdata_out <= ram_w8_l16384_id7_2_1_wdata;
      end else begin
        ram_w8_l16384_id7_2_1_rdata_out <= mem[ram_w8_l16384_id7_2_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l16384_id7_3
(
  input CLK,
  input [12-1:0] ram_w8_l16384_id7_3_0_addr,
  output [8-1:0] ram_w8_l16384_id7_3_0_rdata,
  input [8-1:0] ram_w8_l16384_id7_3_0_wdata,
  input ram_w8_l16384_id7_3_0_wenable,
  input ram_w8_l16384_id7_3_0_enable,
  input [12-1:0] ram_w8_l16384_id7_3_1_addr,
  output [8-1:0] ram_w8_l16384_id7_3_1_rdata,
  input [8-1:0] ram_w8_l16384_id7_3_1_wdata,
  input ram_w8_l16384_id7_3_1_wenable,
  input ram_w8_l16384_id7_3_1_enable
);

  reg [8-1:0] ram_w8_l16384_id7_3_0_rdata_out;
  assign ram_w8_l16384_id7_3_0_rdata = ram_w8_l16384_id7_3_0_rdata_out;
  reg [8-1:0] ram_w8_l16384_id7_3_1_rdata_out;
  assign ram_w8_l16384_id7_3_1_rdata = ram_w8_l16384_id7_3_1_rdata_out;
  reg [8-1:0] mem [0:4096-1];

  always @(posedge CLK) begin
    if(ram_w8_l16384_id7_3_0_enable) begin
      if(ram_w8_l16384_id7_3_0_wenable) begin
        mem[ram_w8_l16384_id7_3_0_addr] <= ram_w8_l16384_id7_3_0_wdata;
        ram_w8_l16384_id7_3_0_rdata_out <= ram_w8_l16384_id7_3_0_wdata;
      end else begin
        ram_w8_l16384_id7_3_0_rdata_out <= mem[ram_w8_l16384_id7_3_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l16384_id7_3_1_enable) begin
      if(ram_w8_l16384_id7_3_1_wenable) begin
        mem[ram_w8_l16384_id7_3_1_addr] <= ram_w8_l16384_id7_3_1_wdata;
        ram_w8_l16384_id7_3_1_rdata_out <= ram_w8_l16384_id7_3_1_wdata;
      end else begin
        ram_w8_l16384_id7_3_1_rdata_out <= mem[ram_w8_l16384_id7_3_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l16384_id8_0
(
  input CLK,
  input [12-1:0] ram_w8_l16384_id8_0_0_addr,
  output [8-1:0] ram_w8_l16384_id8_0_0_rdata,
  input [8-1:0] ram_w8_l16384_id8_0_0_wdata,
  input ram_w8_l16384_id8_0_0_wenable,
  input ram_w8_l16384_id8_0_0_enable,
  input [12-1:0] ram_w8_l16384_id8_0_1_addr,
  output [8-1:0] ram_w8_l16384_id8_0_1_rdata,
  input [8-1:0] ram_w8_l16384_id8_0_1_wdata,
  input ram_w8_l16384_id8_0_1_wenable,
  input ram_w8_l16384_id8_0_1_enable
);

  reg [8-1:0] ram_w8_l16384_id8_0_0_rdata_out;
  assign ram_w8_l16384_id8_0_0_rdata = ram_w8_l16384_id8_0_0_rdata_out;
  reg [8-1:0] ram_w8_l16384_id8_0_1_rdata_out;
  assign ram_w8_l16384_id8_0_1_rdata = ram_w8_l16384_id8_0_1_rdata_out;
  reg [8-1:0] mem [0:4096-1];

  always @(posedge CLK) begin
    if(ram_w8_l16384_id8_0_0_enable) begin
      if(ram_w8_l16384_id8_0_0_wenable) begin
        mem[ram_w8_l16384_id8_0_0_addr] <= ram_w8_l16384_id8_0_0_wdata;
        ram_w8_l16384_id8_0_0_rdata_out <= ram_w8_l16384_id8_0_0_wdata;
      end else begin
        ram_w8_l16384_id8_0_0_rdata_out <= mem[ram_w8_l16384_id8_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l16384_id8_0_1_enable) begin
      if(ram_w8_l16384_id8_0_1_wenable) begin
        mem[ram_w8_l16384_id8_0_1_addr] <= ram_w8_l16384_id8_0_1_wdata;
        ram_w8_l16384_id8_0_1_rdata_out <= ram_w8_l16384_id8_0_1_wdata;
      end else begin
        ram_w8_l16384_id8_0_1_rdata_out <= mem[ram_w8_l16384_id8_0_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l16384_id8_1
(
  input CLK,
  input [12-1:0] ram_w8_l16384_id8_1_0_addr,
  output [8-1:0] ram_w8_l16384_id8_1_0_rdata,
  input [8-1:0] ram_w8_l16384_id8_1_0_wdata,
  input ram_w8_l16384_id8_1_0_wenable,
  input ram_w8_l16384_id8_1_0_enable,
  input [12-1:0] ram_w8_l16384_id8_1_1_addr,
  output [8-1:0] ram_w8_l16384_id8_1_1_rdata,
  input [8-1:0] ram_w8_l16384_id8_1_1_wdata,
  input ram_w8_l16384_id8_1_1_wenable,
  input ram_w8_l16384_id8_1_1_enable
);

  reg [8-1:0] ram_w8_l16384_id8_1_0_rdata_out;
  assign ram_w8_l16384_id8_1_0_rdata = ram_w8_l16384_id8_1_0_rdata_out;
  reg [8-1:0] ram_w8_l16384_id8_1_1_rdata_out;
  assign ram_w8_l16384_id8_1_1_rdata = ram_w8_l16384_id8_1_1_rdata_out;
  reg [8-1:0] mem [0:4096-1];

  always @(posedge CLK) begin
    if(ram_w8_l16384_id8_1_0_enable) begin
      if(ram_w8_l16384_id8_1_0_wenable) begin
        mem[ram_w8_l16384_id8_1_0_addr] <= ram_w8_l16384_id8_1_0_wdata;
        ram_w8_l16384_id8_1_0_rdata_out <= ram_w8_l16384_id8_1_0_wdata;
      end else begin
        ram_w8_l16384_id8_1_0_rdata_out <= mem[ram_w8_l16384_id8_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l16384_id8_1_1_enable) begin
      if(ram_w8_l16384_id8_1_1_wenable) begin
        mem[ram_w8_l16384_id8_1_1_addr] <= ram_w8_l16384_id8_1_1_wdata;
        ram_w8_l16384_id8_1_1_rdata_out <= ram_w8_l16384_id8_1_1_wdata;
      end else begin
        ram_w8_l16384_id8_1_1_rdata_out <= mem[ram_w8_l16384_id8_1_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l16384_id8_2
(
  input CLK,
  input [12-1:0] ram_w8_l16384_id8_2_0_addr,
  output [8-1:0] ram_w8_l16384_id8_2_0_rdata,
  input [8-1:0] ram_w8_l16384_id8_2_0_wdata,
  input ram_w8_l16384_id8_2_0_wenable,
  input ram_w8_l16384_id8_2_0_enable,
  input [12-1:0] ram_w8_l16384_id8_2_1_addr,
  output [8-1:0] ram_w8_l16384_id8_2_1_rdata,
  input [8-1:0] ram_w8_l16384_id8_2_1_wdata,
  input ram_w8_l16384_id8_2_1_wenable,
  input ram_w8_l16384_id8_2_1_enable
);

  reg [8-1:0] ram_w8_l16384_id8_2_0_rdata_out;
  assign ram_w8_l16384_id8_2_0_rdata = ram_w8_l16384_id8_2_0_rdata_out;
  reg [8-1:0] ram_w8_l16384_id8_2_1_rdata_out;
  assign ram_w8_l16384_id8_2_1_rdata = ram_w8_l16384_id8_2_1_rdata_out;
  reg [8-1:0] mem [0:4096-1];

  always @(posedge CLK) begin
    if(ram_w8_l16384_id8_2_0_enable) begin
      if(ram_w8_l16384_id8_2_0_wenable) begin
        mem[ram_w8_l16384_id8_2_0_addr] <= ram_w8_l16384_id8_2_0_wdata;
        ram_w8_l16384_id8_2_0_rdata_out <= ram_w8_l16384_id8_2_0_wdata;
      end else begin
        ram_w8_l16384_id8_2_0_rdata_out <= mem[ram_w8_l16384_id8_2_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l16384_id8_2_1_enable) begin
      if(ram_w8_l16384_id8_2_1_wenable) begin
        mem[ram_w8_l16384_id8_2_1_addr] <= ram_w8_l16384_id8_2_1_wdata;
        ram_w8_l16384_id8_2_1_rdata_out <= ram_w8_l16384_id8_2_1_wdata;
      end else begin
        ram_w8_l16384_id8_2_1_rdata_out <= mem[ram_w8_l16384_id8_2_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l16384_id8_3
(
  input CLK,
  input [12-1:0] ram_w8_l16384_id8_3_0_addr,
  output [8-1:0] ram_w8_l16384_id8_3_0_rdata,
  input [8-1:0] ram_w8_l16384_id8_3_0_wdata,
  input ram_w8_l16384_id8_3_0_wenable,
  input ram_w8_l16384_id8_3_0_enable,
  input [12-1:0] ram_w8_l16384_id8_3_1_addr,
  output [8-1:0] ram_w8_l16384_id8_3_1_rdata,
  input [8-1:0] ram_w8_l16384_id8_3_1_wdata,
  input ram_w8_l16384_id8_3_1_wenable,
  input ram_w8_l16384_id8_3_1_enable
);

  reg [8-1:0] ram_w8_l16384_id8_3_0_rdata_out;
  assign ram_w8_l16384_id8_3_0_rdata = ram_w8_l16384_id8_3_0_rdata_out;
  reg [8-1:0] ram_w8_l16384_id8_3_1_rdata_out;
  assign ram_w8_l16384_id8_3_1_rdata = ram_w8_l16384_id8_3_1_rdata_out;
  reg [8-1:0] mem [0:4096-1];

  always @(posedge CLK) begin
    if(ram_w8_l16384_id8_3_0_enable) begin
      if(ram_w8_l16384_id8_3_0_wenable) begin
        mem[ram_w8_l16384_id8_3_0_addr] <= ram_w8_l16384_id8_3_0_wdata;
        ram_w8_l16384_id8_3_0_rdata_out <= ram_w8_l16384_id8_3_0_wdata;
      end else begin
        ram_w8_l16384_id8_3_0_rdata_out <= mem[ram_w8_l16384_id8_3_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l16384_id8_3_1_enable) begin
      if(ram_w8_l16384_id8_3_1_wenable) begin
        mem[ram_w8_l16384_id8_3_1_addr] <= ram_w8_l16384_id8_3_1_wdata;
        ram_w8_l16384_id8_3_1_rdata_out <= ram_w8_l16384_id8_3_1_wdata;
      end else begin
        ram_w8_l16384_id8_3_1_rdata_out <= mem[ram_w8_l16384_id8_3_1_addr];
      end
    end 
  end


endmodule



module ram_w32_l4096_id0
(
  input CLK,
  input [12-1:0] ram_w32_l4096_id0_0_addr,
  output [32-1:0] ram_w32_l4096_id0_0_rdata,
  input [32-1:0] ram_w32_l4096_id0_0_wdata,
  input ram_w32_l4096_id0_0_wenable,
  input ram_w32_l4096_id0_0_enable,
  input [12-1:0] ram_w32_l4096_id0_1_addr,
  output [32-1:0] ram_w32_l4096_id0_1_rdata,
  input [32-1:0] ram_w32_l4096_id0_1_wdata,
  input ram_w32_l4096_id0_1_wenable,
  input ram_w32_l4096_id0_1_enable
);

  reg [32-1:0] ram_w32_l4096_id0_0_rdata_out;
  assign ram_w32_l4096_id0_0_rdata = ram_w32_l4096_id0_0_rdata_out;
  reg [32-1:0] ram_w32_l4096_id0_1_rdata_out;
  assign ram_w32_l4096_id0_1_rdata = ram_w32_l4096_id0_1_rdata_out;
  reg [32-1:0] mem [0:4096-1];

  always @(posedge CLK) begin
    if(ram_w32_l4096_id0_0_enable) begin
      if(ram_w32_l4096_id0_0_wenable) begin
        mem[ram_w32_l4096_id0_0_addr] <= ram_w32_l4096_id0_0_wdata;
        ram_w32_l4096_id0_0_rdata_out <= ram_w32_l4096_id0_0_wdata;
      end else begin
        ram_w32_l4096_id0_0_rdata_out <= mem[ram_w32_l4096_id0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w32_l4096_id0_1_enable) begin
      if(ram_w32_l4096_id0_1_wenable) begin
        mem[ram_w32_l4096_id0_1_addr] <= ram_w32_l4096_id0_1_wdata;
        ram_w32_l4096_id0_1_rdata_out <= ram_w32_l4096_id0_1_wdata;
      end else begin
        ram_w32_l4096_id0_1_rdata_out <= mem[ram_w32_l4096_id0_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l4096_id0_0
(
  input CLK,
  input [10-1:0] ram_w8_l4096_id0_0_0_addr,
  output [8-1:0] ram_w8_l4096_id0_0_0_rdata,
  input [8-1:0] ram_w8_l4096_id0_0_0_wdata,
  input ram_w8_l4096_id0_0_0_wenable,
  input ram_w8_l4096_id0_0_0_enable,
  input [10-1:0] ram_w8_l4096_id0_0_1_addr,
  output [8-1:0] ram_w8_l4096_id0_0_1_rdata,
  input [8-1:0] ram_w8_l4096_id0_0_1_wdata,
  input ram_w8_l4096_id0_0_1_wenable,
  input ram_w8_l4096_id0_0_1_enable
);

  reg [8-1:0] ram_w8_l4096_id0_0_0_rdata_out;
  assign ram_w8_l4096_id0_0_0_rdata = ram_w8_l4096_id0_0_0_rdata_out;
  reg [8-1:0] ram_w8_l4096_id0_0_1_rdata_out;
  assign ram_w8_l4096_id0_0_1_rdata = ram_w8_l4096_id0_0_1_rdata_out;
  reg [8-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w8_l4096_id0_0_0_enable) begin
      if(ram_w8_l4096_id0_0_0_wenable) begin
        mem[ram_w8_l4096_id0_0_0_addr] <= ram_w8_l4096_id0_0_0_wdata;
        ram_w8_l4096_id0_0_0_rdata_out <= ram_w8_l4096_id0_0_0_wdata;
      end else begin
        ram_w8_l4096_id0_0_0_rdata_out <= mem[ram_w8_l4096_id0_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l4096_id0_0_1_enable) begin
      if(ram_w8_l4096_id0_0_1_wenable) begin
        mem[ram_w8_l4096_id0_0_1_addr] <= ram_w8_l4096_id0_0_1_wdata;
        ram_w8_l4096_id0_0_1_rdata_out <= ram_w8_l4096_id0_0_1_wdata;
      end else begin
        ram_w8_l4096_id0_0_1_rdata_out <= mem[ram_w8_l4096_id0_0_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l4096_id0_1
(
  input CLK,
  input [10-1:0] ram_w8_l4096_id0_1_0_addr,
  output [8-1:0] ram_w8_l4096_id0_1_0_rdata,
  input [8-1:0] ram_w8_l4096_id0_1_0_wdata,
  input ram_w8_l4096_id0_1_0_wenable,
  input ram_w8_l4096_id0_1_0_enable,
  input [10-1:0] ram_w8_l4096_id0_1_1_addr,
  output [8-1:0] ram_w8_l4096_id0_1_1_rdata,
  input [8-1:0] ram_w8_l4096_id0_1_1_wdata,
  input ram_w8_l4096_id0_1_1_wenable,
  input ram_w8_l4096_id0_1_1_enable
);

  reg [8-1:0] ram_w8_l4096_id0_1_0_rdata_out;
  assign ram_w8_l4096_id0_1_0_rdata = ram_w8_l4096_id0_1_0_rdata_out;
  reg [8-1:0] ram_w8_l4096_id0_1_1_rdata_out;
  assign ram_w8_l4096_id0_1_1_rdata = ram_w8_l4096_id0_1_1_rdata_out;
  reg [8-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w8_l4096_id0_1_0_enable) begin
      if(ram_w8_l4096_id0_1_0_wenable) begin
        mem[ram_w8_l4096_id0_1_0_addr] <= ram_w8_l4096_id0_1_0_wdata;
        ram_w8_l4096_id0_1_0_rdata_out <= ram_w8_l4096_id0_1_0_wdata;
      end else begin
        ram_w8_l4096_id0_1_0_rdata_out <= mem[ram_w8_l4096_id0_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l4096_id0_1_1_enable) begin
      if(ram_w8_l4096_id0_1_1_wenable) begin
        mem[ram_w8_l4096_id0_1_1_addr] <= ram_w8_l4096_id0_1_1_wdata;
        ram_w8_l4096_id0_1_1_rdata_out <= ram_w8_l4096_id0_1_1_wdata;
      end else begin
        ram_w8_l4096_id0_1_1_rdata_out <= mem[ram_w8_l4096_id0_1_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l4096_id0_2
(
  input CLK,
  input [10-1:0] ram_w8_l4096_id0_2_0_addr,
  output [8-1:0] ram_w8_l4096_id0_2_0_rdata,
  input [8-1:0] ram_w8_l4096_id0_2_0_wdata,
  input ram_w8_l4096_id0_2_0_wenable,
  input ram_w8_l4096_id0_2_0_enable,
  input [10-1:0] ram_w8_l4096_id0_2_1_addr,
  output [8-1:0] ram_w8_l4096_id0_2_1_rdata,
  input [8-1:0] ram_w8_l4096_id0_2_1_wdata,
  input ram_w8_l4096_id0_2_1_wenable,
  input ram_w8_l4096_id0_2_1_enable
);

  reg [8-1:0] ram_w8_l4096_id0_2_0_rdata_out;
  assign ram_w8_l4096_id0_2_0_rdata = ram_w8_l4096_id0_2_0_rdata_out;
  reg [8-1:0] ram_w8_l4096_id0_2_1_rdata_out;
  assign ram_w8_l4096_id0_2_1_rdata = ram_w8_l4096_id0_2_1_rdata_out;
  reg [8-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w8_l4096_id0_2_0_enable) begin
      if(ram_w8_l4096_id0_2_0_wenable) begin
        mem[ram_w8_l4096_id0_2_0_addr] <= ram_w8_l4096_id0_2_0_wdata;
        ram_w8_l4096_id0_2_0_rdata_out <= ram_w8_l4096_id0_2_0_wdata;
      end else begin
        ram_w8_l4096_id0_2_0_rdata_out <= mem[ram_w8_l4096_id0_2_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l4096_id0_2_1_enable) begin
      if(ram_w8_l4096_id0_2_1_wenable) begin
        mem[ram_w8_l4096_id0_2_1_addr] <= ram_w8_l4096_id0_2_1_wdata;
        ram_w8_l4096_id0_2_1_rdata_out <= ram_w8_l4096_id0_2_1_wdata;
      end else begin
        ram_w8_l4096_id0_2_1_rdata_out <= mem[ram_w8_l4096_id0_2_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l4096_id0_3
(
  input CLK,
  input [10-1:0] ram_w8_l4096_id0_3_0_addr,
  output [8-1:0] ram_w8_l4096_id0_3_0_rdata,
  input [8-1:0] ram_w8_l4096_id0_3_0_wdata,
  input ram_w8_l4096_id0_3_0_wenable,
  input ram_w8_l4096_id0_3_0_enable,
  input [10-1:0] ram_w8_l4096_id0_3_1_addr,
  output [8-1:0] ram_w8_l4096_id0_3_1_rdata,
  input [8-1:0] ram_w8_l4096_id0_3_1_wdata,
  input ram_w8_l4096_id0_3_1_wenable,
  input ram_w8_l4096_id0_3_1_enable
);

  reg [8-1:0] ram_w8_l4096_id0_3_0_rdata_out;
  assign ram_w8_l4096_id0_3_0_rdata = ram_w8_l4096_id0_3_0_rdata_out;
  reg [8-1:0] ram_w8_l4096_id0_3_1_rdata_out;
  assign ram_w8_l4096_id0_3_1_rdata = ram_w8_l4096_id0_3_1_rdata_out;
  reg [8-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w8_l4096_id0_3_0_enable) begin
      if(ram_w8_l4096_id0_3_0_wenable) begin
        mem[ram_w8_l4096_id0_3_0_addr] <= ram_w8_l4096_id0_3_0_wdata;
        ram_w8_l4096_id0_3_0_rdata_out <= ram_w8_l4096_id0_3_0_wdata;
      end else begin
        ram_w8_l4096_id0_3_0_rdata_out <= mem[ram_w8_l4096_id0_3_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l4096_id0_3_1_enable) begin
      if(ram_w8_l4096_id0_3_1_wenable) begin
        mem[ram_w8_l4096_id0_3_1_addr] <= ram_w8_l4096_id0_3_1_wdata;
        ram_w8_l4096_id0_3_1_rdata_out <= ram_w8_l4096_id0_3_1_wdata;
      end else begin
        ram_w8_l4096_id0_3_1_rdata_out <= mem[ram_w8_l4096_id0_3_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l4096_id1_0
(
  input CLK,
  input [10-1:0] ram_w8_l4096_id1_0_0_addr,
  output [8-1:0] ram_w8_l4096_id1_0_0_rdata,
  input [8-1:0] ram_w8_l4096_id1_0_0_wdata,
  input ram_w8_l4096_id1_0_0_wenable,
  input ram_w8_l4096_id1_0_0_enable,
  input [10-1:0] ram_w8_l4096_id1_0_1_addr,
  output [8-1:0] ram_w8_l4096_id1_0_1_rdata,
  input [8-1:0] ram_w8_l4096_id1_0_1_wdata,
  input ram_w8_l4096_id1_0_1_wenable,
  input ram_w8_l4096_id1_0_1_enable
);

  reg [8-1:0] ram_w8_l4096_id1_0_0_rdata_out;
  assign ram_w8_l4096_id1_0_0_rdata = ram_w8_l4096_id1_0_0_rdata_out;
  reg [8-1:0] ram_w8_l4096_id1_0_1_rdata_out;
  assign ram_w8_l4096_id1_0_1_rdata = ram_w8_l4096_id1_0_1_rdata_out;
  reg [8-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w8_l4096_id1_0_0_enable) begin
      if(ram_w8_l4096_id1_0_0_wenable) begin
        mem[ram_w8_l4096_id1_0_0_addr] <= ram_w8_l4096_id1_0_0_wdata;
        ram_w8_l4096_id1_0_0_rdata_out <= ram_w8_l4096_id1_0_0_wdata;
      end else begin
        ram_w8_l4096_id1_0_0_rdata_out <= mem[ram_w8_l4096_id1_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l4096_id1_0_1_enable) begin
      if(ram_w8_l4096_id1_0_1_wenable) begin
        mem[ram_w8_l4096_id1_0_1_addr] <= ram_w8_l4096_id1_0_1_wdata;
        ram_w8_l4096_id1_0_1_rdata_out <= ram_w8_l4096_id1_0_1_wdata;
      end else begin
        ram_w8_l4096_id1_0_1_rdata_out <= mem[ram_w8_l4096_id1_0_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l4096_id1_1
(
  input CLK,
  input [10-1:0] ram_w8_l4096_id1_1_0_addr,
  output [8-1:0] ram_w8_l4096_id1_1_0_rdata,
  input [8-1:0] ram_w8_l4096_id1_1_0_wdata,
  input ram_w8_l4096_id1_1_0_wenable,
  input ram_w8_l4096_id1_1_0_enable,
  input [10-1:0] ram_w8_l4096_id1_1_1_addr,
  output [8-1:0] ram_w8_l4096_id1_1_1_rdata,
  input [8-1:0] ram_w8_l4096_id1_1_1_wdata,
  input ram_w8_l4096_id1_1_1_wenable,
  input ram_w8_l4096_id1_1_1_enable
);

  reg [8-1:0] ram_w8_l4096_id1_1_0_rdata_out;
  assign ram_w8_l4096_id1_1_0_rdata = ram_w8_l4096_id1_1_0_rdata_out;
  reg [8-1:0] ram_w8_l4096_id1_1_1_rdata_out;
  assign ram_w8_l4096_id1_1_1_rdata = ram_w8_l4096_id1_1_1_rdata_out;
  reg [8-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w8_l4096_id1_1_0_enable) begin
      if(ram_w8_l4096_id1_1_0_wenable) begin
        mem[ram_w8_l4096_id1_1_0_addr] <= ram_w8_l4096_id1_1_0_wdata;
        ram_w8_l4096_id1_1_0_rdata_out <= ram_w8_l4096_id1_1_0_wdata;
      end else begin
        ram_w8_l4096_id1_1_0_rdata_out <= mem[ram_w8_l4096_id1_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l4096_id1_1_1_enable) begin
      if(ram_w8_l4096_id1_1_1_wenable) begin
        mem[ram_w8_l4096_id1_1_1_addr] <= ram_w8_l4096_id1_1_1_wdata;
        ram_w8_l4096_id1_1_1_rdata_out <= ram_w8_l4096_id1_1_1_wdata;
      end else begin
        ram_w8_l4096_id1_1_1_rdata_out <= mem[ram_w8_l4096_id1_1_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l4096_id1_2
(
  input CLK,
  input [10-1:0] ram_w8_l4096_id1_2_0_addr,
  output [8-1:0] ram_w8_l4096_id1_2_0_rdata,
  input [8-1:0] ram_w8_l4096_id1_2_0_wdata,
  input ram_w8_l4096_id1_2_0_wenable,
  input ram_w8_l4096_id1_2_0_enable,
  input [10-1:0] ram_w8_l4096_id1_2_1_addr,
  output [8-1:0] ram_w8_l4096_id1_2_1_rdata,
  input [8-1:0] ram_w8_l4096_id1_2_1_wdata,
  input ram_w8_l4096_id1_2_1_wenable,
  input ram_w8_l4096_id1_2_1_enable
);

  reg [8-1:0] ram_w8_l4096_id1_2_0_rdata_out;
  assign ram_w8_l4096_id1_2_0_rdata = ram_w8_l4096_id1_2_0_rdata_out;
  reg [8-1:0] ram_w8_l4096_id1_2_1_rdata_out;
  assign ram_w8_l4096_id1_2_1_rdata = ram_w8_l4096_id1_2_1_rdata_out;
  reg [8-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w8_l4096_id1_2_0_enable) begin
      if(ram_w8_l4096_id1_2_0_wenable) begin
        mem[ram_w8_l4096_id1_2_0_addr] <= ram_w8_l4096_id1_2_0_wdata;
        ram_w8_l4096_id1_2_0_rdata_out <= ram_w8_l4096_id1_2_0_wdata;
      end else begin
        ram_w8_l4096_id1_2_0_rdata_out <= mem[ram_w8_l4096_id1_2_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l4096_id1_2_1_enable) begin
      if(ram_w8_l4096_id1_2_1_wenable) begin
        mem[ram_w8_l4096_id1_2_1_addr] <= ram_w8_l4096_id1_2_1_wdata;
        ram_w8_l4096_id1_2_1_rdata_out <= ram_w8_l4096_id1_2_1_wdata;
      end else begin
        ram_w8_l4096_id1_2_1_rdata_out <= mem[ram_w8_l4096_id1_2_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l4096_id1_3
(
  input CLK,
  input [10-1:0] ram_w8_l4096_id1_3_0_addr,
  output [8-1:0] ram_w8_l4096_id1_3_0_rdata,
  input [8-1:0] ram_w8_l4096_id1_3_0_wdata,
  input ram_w8_l4096_id1_3_0_wenable,
  input ram_w8_l4096_id1_3_0_enable,
  input [10-1:0] ram_w8_l4096_id1_3_1_addr,
  output [8-1:0] ram_w8_l4096_id1_3_1_rdata,
  input [8-1:0] ram_w8_l4096_id1_3_1_wdata,
  input ram_w8_l4096_id1_3_1_wenable,
  input ram_w8_l4096_id1_3_1_enable
);

  reg [8-1:0] ram_w8_l4096_id1_3_0_rdata_out;
  assign ram_w8_l4096_id1_3_0_rdata = ram_w8_l4096_id1_3_0_rdata_out;
  reg [8-1:0] ram_w8_l4096_id1_3_1_rdata_out;
  assign ram_w8_l4096_id1_3_1_rdata = ram_w8_l4096_id1_3_1_rdata_out;
  reg [8-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w8_l4096_id1_3_0_enable) begin
      if(ram_w8_l4096_id1_3_0_wenable) begin
        mem[ram_w8_l4096_id1_3_0_addr] <= ram_w8_l4096_id1_3_0_wdata;
        ram_w8_l4096_id1_3_0_rdata_out <= ram_w8_l4096_id1_3_0_wdata;
      end else begin
        ram_w8_l4096_id1_3_0_rdata_out <= mem[ram_w8_l4096_id1_3_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l4096_id1_3_1_enable) begin
      if(ram_w8_l4096_id1_3_1_wenable) begin
        mem[ram_w8_l4096_id1_3_1_addr] <= ram_w8_l4096_id1_3_1_wdata;
        ram_w8_l4096_id1_3_1_rdata_out <= ram_w8_l4096_id1_3_1_wdata;
      end else begin
        ram_w8_l4096_id1_3_1_rdata_out <= mem[ram_w8_l4096_id1_3_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l4096_id2_0
(
  input CLK,
  input [10-1:0] ram_w8_l4096_id2_0_0_addr,
  output [8-1:0] ram_w8_l4096_id2_0_0_rdata,
  input [8-1:0] ram_w8_l4096_id2_0_0_wdata,
  input ram_w8_l4096_id2_0_0_wenable,
  input ram_w8_l4096_id2_0_0_enable,
  input [10-1:0] ram_w8_l4096_id2_0_1_addr,
  output [8-1:0] ram_w8_l4096_id2_0_1_rdata,
  input [8-1:0] ram_w8_l4096_id2_0_1_wdata,
  input ram_w8_l4096_id2_0_1_wenable,
  input ram_w8_l4096_id2_0_1_enable
);

  reg [8-1:0] ram_w8_l4096_id2_0_0_rdata_out;
  assign ram_w8_l4096_id2_0_0_rdata = ram_w8_l4096_id2_0_0_rdata_out;
  reg [8-1:0] ram_w8_l4096_id2_0_1_rdata_out;
  assign ram_w8_l4096_id2_0_1_rdata = ram_w8_l4096_id2_0_1_rdata_out;
  reg [8-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w8_l4096_id2_0_0_enable) begin
      if(ram_w8_l4096_id2_0_0_wenable) begin
        mem[ram_w8_l4096_id2_0_0_addr] <= ram_w8_l4096_id2_0_0_wdata;
        ram_w8_l4096_id2_0_0_rdata_out <= ram_w8_l4096_id2_0_0_wdata;
      end else begin
        ram_w8_l4096_id2_0_0_rdata_out <= mem[ram_w8_l4096_id2_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l4096_id2_0_1_enable) begin
      if(ram_w8_l4096_id2_0_1_wenable) begin
        mem[ram_w8_l4096_id2_0_1_addr] <= ram_w8_l4096_id2_0_1_wdata;
        ram_w8_l4096_id2_0_1_rdata_out <= ram_w8_l4096_id2_0_1_wdata;
      end else begin
        ram_w8_l4096_id2_0_1_rdata_out <= mem[ram_w8_l4096_id2_0_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l4096_id2_1
(
  input CLK,
  input [10-1:0] ram_w8_l4096_id2_1_0_addr,
  output [8-1:0] ram_w8_l4096_id2_1_0_rdata,
  input [8-1:0] ram_w8_l4096_id2_1_0_wdata,
  input ram_w8_l4096_id2_1_0_wenable,
  input ram_w8_l4096_id2_1_0_enable,
  input [10-1:0] ram_w8_l4096_id2_1_1_addr,
  output [8-1:0] ram_w8_l4096_id2_1_1_rdata,
  input [8-1:0] ram_w8_l4096_id2_1_1_wdata,
  input ram_w8_l4096_id2_1_1_wenable,
  input ram_w8_l4096_id2_1_1_enable
);

  reg [8-1:0] ram_w8_l4096_id2_1_0_rdata_out;
  assign ram_w8_l4096_id2_1_0_rdata = ram_w8_l4096_id2_1_0_rdata_out;
  reg [8-1:0] ram_w8_l4096_id2_1_1_rdata_out;
  assign ram_w8_l4096_id2_1_1_rdata = ram_w8_l4096_id2_1_1_rdata_out;
  reg [8-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w8_l4096_id2_1_0_enable) begin
      if(ram_w8_l4096_id2_1_0_wenable) begin
        mem[ram_w8_l4096_id2_1_0_addr] <= ram_w8_l4096_id2_1_0_wdata;
        ram_w8_l4096_id2_1_0_rdata_out <= ram_w8_l4096_id2_1_0_wdata;
      end else begin
        ram_w8_l4096_id2_1_0_rdata_out <= mem[ram_w8_l4096_id2_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l4096_id2_1_1_enable) begin
      if(ram_w8_l4096_id2_1_1_wenable) begin
        mem[ram_w8_l4096_id2_1_1_addr] <= ram_w8_l4096_id2_1_1_wdata;
        ram_w8_l4096_id2_1_1_rdata_out <= ram_w8_l4096_id2_1_1_wdata;
      end else begin
        ram_w8_l4096_id2_1_1_rdata_out <= mem[ram_w8_l4096_id2_1_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l4096_id2_2
(
  input CLK,
  input [10-1:0] ram_w8_l4096_id2_2_0_addr,
  output [8-1:0] ram_w8_l4096_id2_2_0_rdata,
  input [8-1:0] ram_w8_l4096_id2_2_0_wdata,
  input ram_w8_l4096_id2_2_0_wenable,
  input ram_w8_l4096_id2_2_0_enable,
  input [10-1:0] ram_w8_l4096_id2_2_1_addr,
  output [8-1:0] ram_w8_l4096_id2_2_1_rdata,
  input [8-1:0] ram_w8_l4096_id2_2_1_wdata,
  input ram_w8_l4096_id2_2_1_wenable,
  input ram_w8_l4096_id2_2_1_enable
);

  reg [8-1:0] ram_w8_l4096_id2_2_0_rdata_out;
  assign ram_w8_l4096_id2_2_0_rdata = ram_w8_l4096_id2_2_0_rdata_out;
  reg [8-1:0] ram_w8_l4096_id2_2_1_rdata_out;
  assign ram_w8_l4096_id2_2_1_rdata = ram_w8_l4096_id2_2_1_rdata_out;
  reg [8-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w8_l4096_id2_2_0_enable) begin
      if(ram_w8_l4096_id2_2_0_wenable) begin
        mem[ram_w8_l4096_id2_2_0_addr] <= ram_w8_l4096_id2_2_0_wdata;
        ram_w8_l4096_id2_2_0_rdata_out <= ram_w8_l4096_id2_2_0_wdata;
      end else begin
        ram_w8_l4096_id2_2_0_rdata_out <= mem[ram_w8_l4096_id2_2_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l4096_id2_2_1_enable) begin
      if(ram_w8_l4096_id2_2_1_wenable) begin
        mem[ram_w8_l4096_id2_2_1_addr] <= ram_w8_l4096_id2_2_1_wdata;
        ram_w8_l4096_id2_2_1_rdata_out <= ram_w8_l4096_id2_2_1_wdata;
      end else begin
        ram_w8_l4096_id2_2_1_rdata_out <= mem[ram_w8_l4096_id2_2_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l4096_id2_3
(
  input CLK,
  input [10-1:0] ram_w8_l4096_id2_3_0_addr,
  output [8-1:0] ram_w8_l4096_id2_3_0_rdata,
  input [8-1:0] ram_w8_l4096_id2_3_0_wdata,
  input ram_w8_l4096_id2_3_0_wenable,
  input ram_w8_l4096_id2_3_0_enable,
  input [10-1:0] ram_w8_l4096_id2_3_1_addr,
  output [8-1:0] ram_w8_l4096_id2_3_1_rdata,
  input [8-1:0] ram_w8_l4096_id2_3_1_wdata,
  input ram_w8_l4096_id2_3_1_wenable,
  input ram_w8_l4096_id2_3_1_enable
);

  reg [8-1:0] ram_w8_l4096_id2_3_0_rdata_out;
  assign ram_w8_l4096_id2_3_0_rdata = ram_w8_l4096_id2_3_0_rdata_out;
  reg [8-1:0] ram_w8_l4096_id2_3_1_rdata_out;
  assign ram_w8_l4096_id2_3_1_rdata = ram_w8_l4096_id2_3_1_rdata_out;
  reg [8-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w8_l4096_id2_3_0_enable) begin
      if(ram_w8_l4096_id2_3_0_wenable) begin
        mem[ram_w8_l4096_id2_3_0_addr] <= ram_w8_l4096_id2_3_0_wdata;
        ram_w8_l4096_id2_3_0_rdata_out <= ram_w8_l4096_id2_3_0_wdata;
      end else begin
        ram_w8_l4096_id2_3_0_rdata_out <= mem[ram_w8_l4096_id2_3_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l4096_id2_3_1_enable) begin
      if(ram_w8_l4096_id2_3_1_wenable) begin
        mem[ram_w8_l4096_id2_3_1_addr] <= ram_w8_l4096_id2_3_1_wdata;
        ram_w8_l4096_id2_3_1_rdata_out <= ram_w8_l4096_id2_3_1_wdata;
      end else begin
        ram_w8_l4096_id2_3_1_rdata_out <= mem[ram_w8_l4096_id2_3_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l4096_id3_0
(
  input CLK,
  input [10-1:0] ram_w8_l4096_id3_0_0_addr,
  output [8-1:0] ram_w8_l4096_id3_0_0_rdata,
  input [8-1:0] ram_w8_l4096_id3_0_0_wdata,
  input ram_w8_l4096_id3_0_0_wenable,
  input ram_w8_l4096_id3_0_0_enable,
  input [10-1:0] ram_w8_l4096_id3_0_1_addr,
  output [8-1:0] ram_w8_l4096_id3_0_1_rdata,
  input [8-1:0] ram_w8_l4096_id3_0_1_wdata,
  input ram_w8_l4096_id3_0_1_wenable,
  input ram_w8_l4096_id3_0_1_enable
);

  reg [8-1:0] ram_w8_l4096_id3_0_0_rdata_out;
  assign ram_w8_l4096_id3_0_0_rdata = ram_w8_l4096_id3_0_0_rdata_out;
  reg [8-1:0] ram_w8_l4096_id3_0_1_rdata_out;
  assign ram_w8_l4096_id3_0_1_rdata = ram_w8_l4096_id3_0_1_rdata_out;
  reg [8-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w8_l4096_id3_0_0_enable) begin
      if(ram_w8_l4096_id3_0_0_wenable) begin
        mem[ram_w8_l4096_id3_0_0_addr] <= ram_w8_l4096_id3_0_0_wdata;
        ram_w8_l4096_id3_0_0_rdata_out <= ram_w8_l4096_id3_0_0_wdata;
      end else begin
        ram_w8_l4096_id3_0_0_rdata_out <= mem[ram_w8_l4096_id3_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l4096_id3_0_1_enable) begin
      if(ram_w8_l4096_id3_0_1_wenable) begin
        mem[ram_w8_l4096_id3_0_1_addr] <= ram_w8_l4096_id3_0_1_wdata;
        ram_w8_l4096_id3_0_1_rdata_out <= ram_w8_l4096_id3_0_1_wdata;
      end else begin
        ram_w8_l4096_id3_0_1_rdata_out <= mem[ram_w8_l4096_id3_0_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l4096_id3_1
(
  input CLK,
  input [10-1:0] ram_w8_l4096_id3_1_0_addr,
  output [8-1:0] ram_w8_l4096_id3_1_0_rdata,
  input [8-1:0] ram_w8_l4096_id3_1_0_wdata,
  input ram_w8_l4096_id3_1_0_wenable,
  input ram_w8_l4096_id3_1_0_enable,
  input [10-1:0] ram_w8_l4096_id3_1_1_addr,
  output [8-1:0] ram_w8_l4096_id3_1_1_rdata,
  input [8-1:0] ram_w8_l4096_id3_1_1_wdata,
  input ram_w8_l4096_id3_1_1_wenable,
  input ram_w8_l4096_id3_1_1_enable
);

  reg [8-1:0] ram_w8_l4096_id3_1_0_rdata_out;
  assign ram_w8_l4096_id3_1_0_rdata = ram_w8_l4096_id3_1_0_rdata_out;
  reg [8-1:0] ram_w8_l4096_id3_1_1_rdata_out;
  assign ram_w8_l4096_id3_1_1_rdata = ram_w8_l4096_id3_1_1_rdata_out;
  reg [8-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w8_l4096_id3_1_0_enable) begin
      if(ram_w8_l4096_id3_1_0_wenable) begin
        mem[ram_w8_l4096_id3_1_0_addr] <= ram_w8_l4096_id3_1_0_wdata;
        ram_w8_l4096_id3_1_0_rdata_out <= ram_w8_l4096_id3_1_0_wdata;
      end else begin
        ram_w8_l4096_id3_1_0_rdata_out <= mem[ram_w8_l4096_id3_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l4096_id3_1_1_enable) begin
      if(ram_w8_l4096_id3_1_1_wenable) begin
        mem[ram_w8_l4096_id3_1_1_addr] <= ram_w8_l4096_id3_1_1_wdata;
        ram_w8_l4096_id3_1_1_rdata_out <= ram_w8_l4096_id3_1_1_wdata;
      end else begin
        ram_w8_l4096_id3_1_1_rdata_out <= mem[ram_w8_l4096_id3_1_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l4096_id3_2
(
  input CLK,
  input [10-1:0] ram_w8_l4096_id3_2_0_addr,
  output [8-1:0] ram_w8_l4096_id3_2_0_rdata,
  input [8-1:0] ram_w8_l4096_id3_2_0_wdata,
  input ram_w8_l4096_id3_2_0_wenable,
  input ram_w8_l4096_id3_2_0_enable,
  input [10-1:0] ram_w8_l4096_id3_2_1_addr,
  output [8-1:0] ram_w8_l4096_id3_2_1_rdata,
  input [8-1:0] ram_w8_l4096_id3_2_1_wdata,
  input ram_w8_l4096_id3_2_1_wenable,
  input ram_w8_l4096_id3_2_1_enable
);

  reg [8-1:0] ram_w8_l4096_id3_2_0_rdata_out;
  assign ram_w8_l4096_id3_2_0_rdata = ram_w8_l4096_id3_2_0_rdata_out;
  reg [8-1:0] ram_w8_l4096_id3_2_1_rdata_out;
  assign ram_w8_l4096_id3_2_1_rdata = ram_w8_l4096_id3_2_1_rdata_out;
  reg [8-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w8_l4096_id3_2_0_enable) begin
      if(ram_w8_l4096_id3_2_0_wenable) begin
        mem[ram_w8_l4096_id3_2_0_addr] <= ram_w8_l4096_id3_2_0_wdata;
        ram_w8_l4096_id3_2_0_rdata_out <= ram_w8_l4096_id3_2_0_wdata;
      end else begin
        ram_w8_l4096_id3_2_0_rdata_out <= mem[ram_w8_l4096_id3_2_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l4096_id3_2_1_enable) begin
      if(ram_w8_l4096_id3_2_1_wenable) begin
        mem[ram_w8_l4096_id3_2_1_addr] <= ram_w8_l4096_id3_2_1_wdata;
        ram_w8_l4096_id3_2_1_rdata_out <= ram_w8_l4096_id3_2_1_wdata;
      end else begin
        ram_w8_l4096_id3_2_1_rdata_out <= mem[ram_w8_l4096_id3_2_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l4096_id3_3
(
  input CLK,
  input [10-1:0] ram_w8_l4096_id3_3_0_addr,
  output [8-1:0] ram_w8_l4096_id3_3_0_rdata,
  input [8-1:0] ram_w8_l4096_id3_3_0_wdata,
  input ram_w8_l4096_id3_3_0_wenable,
  input ram_w8_l4096_id3_3_0_enable,
  input [10-1:0] ram_w8_l4096_id3_3_1_addr,
  output [8-1:0] ram_w8_l4096_id3_3_1_rdata,
  input [8-1:0] ram_w8_l4096_id3_3_1_wdata,
  input ram_w8_l4096_id3_3_1_wenable,
  input ram_w8_l4096_id3_3_1_enable
);

  reg [8-1:0] ram_w8_l4096_id3_3_0_rdata_out;
  assign ram_w8_l4096_id3_3_0_rdata = ram_w8_l4096_id3_3_0_rdata_out;
  reg [8-1:0] ram_w8_l4096_id3_3_1_rdata_out;
  assign ram_w8_l4096_id3_3_1_rdata = ram_w8_l4096_id3_3_1_rdata_out;
  reg [8-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w8_l4096_id3_3_0_enable) begin
      if(ram_w8_l4096_id3_3_0_wenable) begin
        mem[ram_w8_l4096_id3_3_0_addr] <= ram_w8_l4096_id3_3_0_wdata;
        ram_w8_l4096_id3_3_0_rdata_out <= ram_w8_l4096_id3_3_0_wdata;
      end else begin
        ram_w8_l4096_id3_3_0_rdata_out <= mem[ram_w8_l4096_id3_3_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l4096_id3_3_1_enable) begin
      if(ram_w8_l4096_id3_3_1_wenable) begin
        mem[ram_w8_l4096_id3_3_1_addr] <= ram_w8_l4096_id3_3_1_wdata;
        ram_w8_l4096_id3_3_1_rdata_out <= ram_w8_l4096_id3_3_1_wdata;
      end else begin
        ram_w8_l4096_id3_3_1_rdata_out <= mem[ram_w8_l4096_id3_3_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l4096_id4_0
(
  input CLK,
  input [10-1:0] ram_w8_l4096_id4_0_0_addr,
  output [8-1:0] ram_w8_l4096_id4_0_0_rdata,
  input [8-1:0] ram_w8_l4096_id4_0_0_wdata,
  input ram_w8_l4096_id4_0_0_wenable,
  input ram_w8_l4096_id4_0_0_enable,
  input [10-1:0] ram_w8_l4096_id4_0_1_addr,
  output [8-1:0] ram_w8_l4096_id4_0_1_rdata,
  input [8-1:0] ram_w8_l4096_id4_0_1_wdata,
  input ram_w8_l4096_id4_0_1_wenable,
  input ram_w8_l4096_id4_0_1_enable
);

  reg [8-1:0] ram_w8_l4096_id4_0_0_rdata_out;
  assign ram_w8_l4096_id4_0_0_rdata = ram_w8_l4096_id4_0_0_rdata_out;
  reg [8-1:0] ram_w8_l4096_id4_0_1_rdata_out;
  assign ram_w8_l4096_id4_0_1_rdata = ram_w8_l4096_id4_0_1_rdata_out;
  reg [8-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w8_l4096_id4_0_0_enable) begin
      if(ram_w8_l4096_id4_0_0_wenable) begin
        mem[ram_w8_l4096_id4_0_0_addr] <= ram_w8_l4096_id4_0_0_wdata;
        ram_w8_l4096_id4_0_0_rdata_out <= ram_w8_l4096_id4_0_0_wdata;
      end else begin
        ram_w8_l4096_id4_0_0_rdata_out <= mem[ram_w8_l4096_id4_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l4096_id4_0_1_enable) begin
      if(ram_w8_l4096_id4_0_1_wenable) begin
        mem[ram_w8_l4096_id4_0_1_addr] <= ram_w8_l4096_id4_0_1_wdata;
        ram_w8_l4096_id4_0_1_rdata_out <= ram_w8_l4096_id4_0_1_wdata;
      end else begin
        ram_w8_l4096_id4_0_1_rdata_out <= mem[ram_w8_l4096_id4_0_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l4096_id4_1
(
  input CLK,
  input [10-1:0] ram_w8_l4096_id4_1_0_addr,
  output [8-1:0] ram_w8_l4096_id4_1_0_rdata,
  input [8-1:0] ram_w8_l4096_id4_1_0_wdata,
  input ram_w8_l4096_id4_1_0_wenable,
  input ram_w8_l4096_id4_1_0_enable,
  input [10-1:0] ram_w8_l4096_id4_1_1_addr,
  output [8-1:0] ram_w8_l4096_id4_1_1_rdata,
  input [8-1:0] ram_w8_l4096_id4_1_1_wdata,
  input ram_w8_l4096_id4_1_1_wenable,
  input ram_w8_l4096_id4_1_1_enable
);

  reg [8-1:0] ram_w8_l4096_id4_1_0_rdata_out;
  assign ram_w8_l4096_id4_1_0_rdata = ram_w8_l4096_id4_1_0_rdata_out;
  reg [8-1:0] ram_w8_l4096_id4_1_1_rdata_out;
  assign ram_w8_l4096_id4_1_1_rdata = ram_w8_l4096_id4_1_1_rdata_out;
  reg [8-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w8_l4096_id4_1_0_enable) begin
      if(ram_w8_l4096_id4_1_0_wenable) begin
        mem[ram_w8_l4096_id4_1_0_addr] <= ram_w8_l4096_id4_1_0_wdata;
        ram_w8_l4096_id4_1_0_rdata_out <= ram_w8_l4096_id4_1_0_wdata;
      end else begin
        ram_w8_l4096_id4_1_0_rdata_out <= mem[ram_w8_l4096_id4_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l4096_id4_1_1_enable) begin
      if(ram_w8_l4096_id4_1_1_wenable) begin
        mem[ram_w8_l4096_id4_1_1_addr] <= ram_w8_l4096_id4_1_1_wdata;
        ram_w8_l4096_id4_1_1_rdata_out <= ram_w8_l4096_id4_1_1_wdata;
      end else begin
        ram_w8_l4096_id4_1_1_rdata_out <= mem[ram_w8_l4096_id4_1_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l4096_id4_2
(
  input CLK,
  input [10-1:0] ram_w8_l4096_id4_2_0_addr,
  output [8-1:0] ram_w8_l4096_id4_2_0_rdata,
  input [8-1:0] ram_w8_l4096_id4_2_0_wdata,
  input ram_w8_l4096_id4_2_0_wenable,
  input ram_w8_l4096_id4_2_0_enable,
  input [10-1:0] ram_w8_l4096_id4_2_1_addr,
  output [8-1:0] ram_w8_l4096_id4_2_1_rdata,
  input [8-1:0] ram_w8_l4096_id4_2_1_wdata,
  input ram_w8_l4096_id4_2_1_wenable,
  input ram_w8_l4096_id4_2_1_enable
);

  reg [8-1:0] ram_w8_l4096_id4_2_0_rdata_out;
  assign ram_w8_l4096_id4_2_0_rdata = ram_w8_l4096_id4_2_0_rdata_out;
  reg [8-1:0] ram_w8_l4096_id4_2_1_rdata_out;
  assign ram_w8_l4096_id4_2_1_rdata = ram_w8_l4096_id4_2_1_rdata_out;
  reg [8-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w8_l4096_id4_2_0_enable) begin
      if(ram_w8_l4096_id4_2_0_wenable) begin
        mem[ram_w8_l4096_id4_2_0_addr] <= ram_w8_l4096_id4_2_0_wdata;
        ram_w8_l4096_id4_2_0_rdata_out <= ram_w8_l4096_id4_2_0_wdata;
      end else begin
        ram_w8_l4096_id4_2_0_rdata_out <= mem[ram_w8_l4096_id4_2_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l4096_id4_2_1_enable) begin
      if(ram_w8_l4096_id4_2_1_wenable) begin
        mem[ram_w8_l4096_id4_2_1_addr] <= ram_w8_l4096_id4_2_1_wdata;
        ram_w8_l4096_id4_2_1_rdata_out <= ram_w8_l4096_id4_2_1_wdata;
      end else begin
        ram_w8_l4096_id4_2_1_rdata_out <= mem[ram_w8_l4096_id4_2_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l4096_id4_3
(
  input CLK,
  input [10-1:0] ram_w8_l4096_id4_3_0_addr,
  output [8-1:0] ram_w8_l4096_id4_3_0_rdata,
  input [8-1:0] ram_w8_l4096_id4_3_0_wdata,
  input ram_w8_l4096_id4_3_0_wenable,
  input ram_w8_l4096_id4_3_0_enable,
  input [10-1:0] ram_w8_l4096_id4_3_1_addr,
  output [8-1:0] ram_w8_l4096_id4_3_1_rdata,
  input [8-1:0] ram_w8_l4096_id4_3_1_wdata,
  input ram_w8_l4096_id4_3_1_wenable,
  input ram_w8_l4096_id4_3_1_enable
);

  reg [8-1:0] ram_w8_l4096_id4_3_0_rdata_out;
  assign ram_w8_l4096_id4_3_0_rdata = ram_w8_l4096_id4_3_0_rdata_out;
  reg [8-1:0] ram_w8_l4096_id4_3_1_rdata_out;
  assign ram_w8_l4096_id4_3_1_rdata = ram_w8_l4096_id4_3_1_rdata_out;
  reg [8-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w8_l4096_id4_3_0_enable) begin
      if(ram_w8_l4096_id4_3_0_wenable) begin
        mem[ram_w8_l4096_id4_3_0_addr] <= ram_w8_l4096_id4_3_0_wdata;
        ram_w8_l4096_id4_3_0_rdata_out <= ram_w8_l4096_id4_3_0_wdata;
      end else begin
        ram_w8_l4096_id4_3_0_rdata_out <= mem[ram_w8_l4096_id4_3_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l4096_id4_3_1_enable) begin
      if(ram_w8_l4096_id4_3_1_wenable) begin
        mem[ram_w8_l4096_id4_3_1_addr] <= ram_w8_l4096_id4_3_1_wdata;
        ram_w8_l4096_id4_3_1_rdata_out <= ram_w8_l4096_id4_3_1_wdata;
      end else begin
        ram_w8_l4096_id4_3_1_rdata_out <= mem[ram_w8_l4096_id4_3_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l4096_id5_0
(
  input CLK,
  input [10-1:0] ram_w8_l4096_id5_0_0_addr,
  output [8-1:0] ram_w8_l4096_id5_0_0_rdata,
  input [8-1:0] ram_w8_l4096_id5_0_0_wdata,
  input ram_w8_l4096_id5_0_0_wenable,
  input ram_w8_l4096_id5_0_0_enable,
  input [10-1:0] ram_w8_l4096_id5_0_1_addr,
  output [8-1:0] ram_w8_l4096_id5_0_1_rdata,
  input [8-1:0] ram_w8_l4096_id5_0_1_wdata,
  input ram_w8_l4096_id5_0_1_wenable,
  input ram_w8_l4096_id5_0_1_enable
);

  reg [8-1:0] ram_w8_l4096_id5_0_0_rdata_out;
  assign ram_w8_l4096_id5_0_0_rdata = ram_w8_l4096_id5_0_0_rdata_out;
  reg [8-1:0] ram_w8_l4096_id5_0_1_rdata_out;
  assign ram_w8_l4096_id5_0_1_rdata = ram_w8_l4096_id5_0_1_rdata_out;
  reg [8-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w8_l4096_id5_0_0_enable) begin
      if(ram_w8_l4096_id5_0_0_wenable) begin
        mem[ram_w8_l4096_id5_0_0_addr] <= ram_w8_l4096_id5_0_0_wdata;
        ram_w8_l4096_id5_0_0_rdata_out <= ram_w8_l4096_id5_0_0_wdata;
      end else begin
        ram_w8_l4096_id5_0_0_rdata_out <= mem[ram_w8_l4096_id5_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l4096_id5_0_1_enable) begin
      if(ram_w8_l4096_id5_0_1_wenable) begin
        mem[ram_w8_l4096_id5_0_1_addr] <= ram_w8_l4096_id5_0_1_wdata;
        ram_w8_l4096_id5_0_1_rdata_out <= ram_w8_l4096_id5_0_1_wdata;
      end else begin
        ram_w8_l4096_id5_0_1_rdata_out <= mem[ram_w8_l4096_id5_0_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l4096_id5_1
(
  input CLK,
  input [10-1:0] ram_w8_l4096_id5_1_0_addr,
  output [8-1:0] ram_w8_l4096_id5_1_0_rdata,
  input [8-1:0] ram_w8_l4096_id5_1_0_wdata,
  input ram_w8_l4096_id5_1_0_wenable,
  input ram_w8_l4096_id5_1_0_enable,
  input [10-1:0] ram_w8_l4096_id5_1_1_addr,
  output [8-1:0] ram_w8_l4096_id5_1_1_rdata,
  input [8-1:0] ram_w8_l4096_id5_1_1_wdata,
  input ram_w8_l4096_id5_1_1_wenable,
  input ram_w8_l4096_id5_1_1_enable
);

  reg [8-1:0] ram_w8_l4096_id5_1_0_rdata_out;
  assign ram_w8_l4096_id5_1_0_rdata = ram_w8_l4096_id5_1_0_rdata_out;
  reg [8-1:0] ram_w8_l4096_id5_1_1_rdata_out;
  assign ram_w8_l4096_id5_1_1_rdata = ram_w8_l4096_id5_1_1_rdata_out;
  reg [8-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w8_l4096_id5_1_0_enable) begin
      if(ram_w8_l4096_id5_1_0_wenable) begin
        mem[ram_w8_l4096_id5_1_0_addr] <= ram_w8_l4096_id5_1_0_wdata;
        ram_w8_l4096_id5_1_0_rdata_out <= ram_w8_l4096_id5_1_0_wdata;
      end else begin
        ram_w8_l4096_id5_1_0_rdata_out <= mem[ram_w8_l4096_id5_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l4096_id5_1_1_enable) begin
      if(ram_w8_l4096_id5_1_1_wenable) begin
        mem[ram_w8_l4096_id5_1_1_addr] <= ram_w8_l4096_id5_1_1_wdata;
        ram_w8_l4096_id5_1_1_rdata_out <= ram_w8_l4096_id5_1_1_wdata;
      end else begin
        ram_w8_l4096_id5_1_1_rdata_out <= mem[ram_w8_l4096_id5_1_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l4096_id5_2
(
  input CLK,
  input [10-1:0] ram_w8_l4096_id5_2_0_addr,
  output [8-1:0] ram_w8_l4096_id5_2_0_rdata,
  input [8-1:0] ram_w8_l4096_id5_2_0_wdata,
  input ram_w8_l4096_id5_2_0_wenable,
  input ram_w8_l4096_id5_2_0_enable,
  input [10-1:0] ram_w8_l4096_id5_2_1_addr,
  output [8-1:0] ram_w8_l4096_id5_2_1_rdata,
  input [8-1:0] ram_w8_l4096_id5_2_1_wdata,
  input ram_w8_l4096_id5_2_1_wenable,
  input ram_w8_l4096_id5_2_1_enable
);

  reg [8-1:0] ram_w8_l4096_id5_2_0_rdata_out;
  assign ram_w8_l4096_id5_2_0_rdata = ram_w8_l4096_id5_2_0_rdata_out;
  reg [8-1:0] ram_w8_l4096_id5_2_1_rdata_out;
  assign ram_w8_l4096_id5_2_1_rdata = ram_w8_l4096_id5_2_1_rdata_out;
  reg [8-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w8_l4096_id5_2_0_enable) begin
      if(ram_w8_l4096_id5_2_0_wenable) begin
        mem[ram_w8_l4096_id5_2_0_addr] <= ram_w8_l4096_id5_2_0_wdata;
        ram_w8_l4096_id5_2_0_rdata_out <= ram_w8_l4096_id5_2_0_wdata;
      end else begin
        ram_w8_l4096_id5_2_0_rdata_out <= mem[ram_w8_l4096_id5_2_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l4096_id5_2_1_enable) begin
      if(ram_w8_l4096_id5_2_1_wenable) begin
        mem[ram_w8_l4096_id5_2_1_addr] <= ram_w8_l4096_id5_2_1_wdata;
        ram_w8_l4096_id5_2_1_rdata_out <= ram_w8_l4096_id5_2_1_wdata;
      end else begin
        ram_w8_l4096_id5_2_1_rdata_out <= mem[ram_w8_l4096_id5_2_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l4096_id5_3
(
  input CLK,
  input [10-1:0] ram_w8_l4096_id5_3_0_addr,
  output [8-1:0] ram_w8_l4096_id5_3_0_rdata,
  input [8-1:0] ram_w8_l4096_id5_3_0_wdata,
  input ram_w8_l4096_id5_3_0_wenable,
  input ram_w8_l4096_id5_3_0_enable,
  input [10-1:0] ram_w8_l4096_id5_3_1_addr,
  output [8-1:0] ram_w8_l4096_id5_3_1_rdata,
  input [8-1:0] ram_w8_l4096_id5_3_1_wdata,
  input ram_w8_l4096_id5_3_1_wenable,
  input ram_w8_l4096_id5_3_1_enable
);

  reg [8-1:0] ram_w8_l4096_id5_3_0_rdata_out;
  assign ram_w8_l4096_id5_3_0_rdata = ram_w8_l4096_id5_3_0_rdata_out;
  reg [8-1:0] ram_w8_l4096_id5_3_1_rdata_out;
  assign ram_w8_l4096_id5_3_1_rdata = ram_w8_l4096_id5_3_1_rdata_out;
  reg [8-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w8_l4096_id5_3_0_enable) begin
      if(ram_w8_l4096_id5_3_0_wenable) begin
        mem[ram_w8_l4096_id5_3_0_addr] <= ram_w8_l4096_id5_3_0_wdata;
        ram_w8_l4096_id5_3_0_rdata_out <= ram_w8_l4096_id5_3_0_wdata;
      end else begin
        ram_w8_l4096_id5_3_0_rdata_out <= mem[ram_w8_l4096_id5_3_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l4096_id5_3_1_enable) begin
      if(ram_w8_l4096_id5_3_1_wenable) begin
        mem[ram_w8_l4096_id5_3_1_addr] <= ram_w8_l4096_id5_3_1_wdata;
        ram_w8_l4096_id5_3_1_rdata_out <= ram_w8_l4096_id5_3_1_wdata;
      end else begin
        ram_w8_l4096_id5_3_1_rdata_out <= mem[ram_w8_l4096_id5_3_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l4096_id6_0
(
  input CLK,
  input [10-1:0] ram_w8_l4096_id6_0_0_addr,
  output [8-1:0] ram_w8_l4096_id6_0_0_rdata,
  input [8-1:0] ram_w8_l4096_id6_0_0_wdata,
  input ram_w8_l4096_id6_0_0_wenable,
  input ram_w8_l4096_id6_0_0_enable,
  input [10-1:0] ram_w8_l4096_id6_0_1_addr,
  output [8-1:0] ram_w8_l4096_id6_0_1_rdata,
  input [8-1:0] ram_w8_l4096_id6_0_1_wdata,
  input ram_w8_l4096_id6_0_1_wenable,
  input ram_w8_l4096_id6_0_1_enable
);

  reg [8-1:0] ram_w8_l4096_id6_0_0_rdata_out;
  assign ram_w8_l4096_id6_0_0_rdata = ram_w8_l4096_id6_0_0_rdata_out;
  reg [8-1:0] ram_w8_l4096_id6_0_1_rdata_out;
  assign ram_w8_l4096_id6_0_1_rdata = ram_w8_l4096_id6_0_1_rdata_out;
  reg [8-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w8_l4096_id6_0_0_enable) begin
      if(ram_w8_l4096_id6_0_0_wenable) begin
        mem[ram_w8_l4096_id6_0_0_addr] <= ram_w8_l4096_id6_0_0_wdata;
        ram_w8_l4096_id6_0_0_rdata_out <= ram_w8_l4096_id6_0_0_wdata;
      end else begin
        ram_w8_l4096_id6_0_0_rdata_out <= mem[ram_w8_l4096_id6_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l4096_id6_0_1_enable) begin
      if(ram_w8_l4096_id6_0_1_wenable) begin
        mem[ram_w8_l4096_id6_0_1_addr] <= ram_w8_l4096_id6_0_1_wdata;
        ram_w8_l4096_id6_0_1_rdata_out <= ram_w8_l4096_id6_0_1_wdata;
      end else begin
        ram_w8_l4096_id6_0_1_rdata_out <= mem[ram_w8_l4096_id6_0_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l4096_id6_1
(
  input CLK,
  input [10-1:0] ram_w8_l4096_id6_1_0_addr,
  output [8-1:0] ram_w8_l4096_id6_1_0_rdata,
  input [8-1:0] ram_w8_l4096_id6_1_0_wdata,
  input ram_w8_l4096_id6_1_0_wenable,
  input ram_w8_l4096_id6_1_0_enable,
  input [10-1:0] ram_w8_l4096_id6_1_1_addr,
  output [8-1:0] ram_w8_l4096_id6_1_1_rdata,
  input [8-1:0] ram_w8_l4096_id6_1_1_wdata,
  input ram_w8_l4096_id6_1_1_wenable,
  input ram_w8_l4096_id6_1_1_enable
);

  reg [8-1:0] ram_w8_l4096_id6_1_0_rdata_out;
  assign ram_w8_l4096_id6_1_0_rdata = ram_w8_l4096_id6_1_0_rdata_out;
  reg [8-1:0] ram_w8_l4096_id6_1_1_rdata_out;
  assign ram_w8_l4096_id6_1_1_rdata = ram_w8_l4096_id6_1_1_rdata_out;
  reg [8-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w8_l4096_id6_1_0_enable) begin
      if(ram_w8_l4096_id6_1_0_wenable) begin
        mem[ram_w8_l4096_id6_1_0_addr] <= ram_w8_l4096_id6_1_0_wdata;
        ram_w8_l4096_id6_1_0_rdata_out <= ram_w8_l4096_id6_1_0_wdata;
      end else begin
        ram_w8_l4096_id6_1_0_rdata_out <= mem[ram_w8_l4096_id6_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l4096_id6_1_1_enable) begin
      if(ram_w8_l4096_id6_1_1_wenable) begin
        mem[ram_w8_l4096_id6_1_1_addr] <= ram_w8_l4096_id6_1_1_wdata;
        ram_w8_l4096_id6_1_1_rdata_out <= ram_w8_l4096_id6_1_1_wdata;
      end else begin
        ram_w8_l4096_id6_1_1_rdata_out <= mem[ram_w8_l4096_id6_1_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l4096_id6_2
(
  input CLK,
  input [10-1:0] ram_w8_l4096_id6_2_0_addr,
  output [8-1:0] ram_w8_l4096_id6_2_0_rdata,
  input [8-1:0] ram_w8_l4096_id6_2_0_wdata,
  input ram_w8_l4096_id6_2_0_wenable,
  input ram_w8_l4096_id6_2_0_enable,
  input [10-1:0] ram_w8_l4096_id6_2_1_addr,
  output [8-1:0] ram_w8_l4096_id6_2_1_rdata,
  input [8-1:0] ram_w8_l4096_id6_2_1_wdata,
  input ram_w8_l4096_id6_2_1_wenable,
  input ram_w8_l4096_id6_2_1_enable
);

  reg [8-1:0] ram_w8_l4096_id6_2_0_rdata_out;
  assign ram_w8_l4096_id6_2_0_rdata = ram_w8_l4096_id6_2_0_rdata_out;
  reg [8-1:0] ram_w8_l4096_id6_2_1_rdata_out;
  assign ram_w8_l4096_id6_2_1_rdata = ram_w8_l4096_id6_2_1_rdata_out;
  reg [8-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w8_l4096_id6_2_0_enable) begin
      if(ram_w8_l4096_id6_2_0_wenable) begin
        mem[ram_w8_l4096_id6_2_0_addr] <= ram_w8_l4096_id6_2_0_wdata;
        ram_w8_l4096_id6_2_0_rdata_out <= ram_w8_l4096_id6_2_0_wdata;
      end else begin
        ram_w8_l4096_id6_2_0_rdata_out <= mem[ram_w8_l4096_id6_2_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l4096_id6_2_1_enable) begin
      if(ram_w8_l4096_id6_2_1_wenable) begin
        mem[ram_w8_l4096_id6_2_1_addr] <= ram_w8_l4096_id6_2_1_wdata;
        ram_w8_l4096_id6_2_1_rdata_out <= ram_w8_l4096_id6_2_1_wdata;
      end else begin
        ram_w8_l4096_id6_2_1_rdata_out <= mem[ram_w8_l4096_id6_2_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l4096_id6_3
(
  input CLK,
  input [10-1:0] ram_w8_l4096_id6_3_0_addr,
  output [8-1:0] ram_w8_l4096_id6_3_0_rdata,
  input [8-1:0] ram_w8_l4096_id6_3_0_wdata,
  input ram_w8_l4096_id6_3_0_wenable,
  input ram_w8_l4096_id6_3_0_enable,
  input [10-1:0] ram_w8_l4096_id6_3_1_addr,
  output [8-1:0] ram_w8_l4096_id6_3_1_rdata,
  input [8-1:0] ram_w8_l4096_id6_3_1_wdata,
  input ram_w8_l4096_id6_3_1_wenable,
  input ram_w8_l4096_id6_3_1_enable
);

  reg [8-1:0] ram_w8_l4096_id6_3_0_rdata_out;
  assign ram_w8_l4096_id6_3_0_rdata = ram_w8_l4096_id6_3_0_rdata_out;
  reg [8-1:0] ram_w8_l4096_id6_3_1_rdata_out;
  assign ram_w8_l4096_id6_3_1_rdata = ram_w8_l4096_id6_3_1_rdata_out;
  reg [8-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w8_l4096_id6_3_0_enable) begin
      if(ram_w8_l4096_id6_3_0_wenable) begin
        mem[ram_w8_l4096_id6_3_0_addr] <= ram_w8_l4096_id6_3_0_wdata;
        ram_w8_l4096_id6_3_0_rdata_out <= ram_w8_l4096_id6_3_0_wdata;
      end else begin
        ram_w8_l4096_id6_3_0_rdata_out <= mem[ram_w8_l4096_id6_3_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l4096_id6_3_1_enable) begin
      if(ram_w8_l4096_id6_3_1_wenable) begin
        mem[ram_w8_l4096_id6_3_1_addr] <= ram_w8_l4096_id6_3_1_wdata;
        ram_w8_l4096_id6_3_1_rdata_out <= ram_w8_l4096_id6_3_1_wdata;
      end else begin
        ram_w8_l4096_id6_3_1_rdata_out <= mem[ram_w8_l4096_id6_3_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l4096_id7_0
(
  input CLK,
  input [10-1:0] ram_w8_l4096_id7_0_0_addr,
  output [8-1:0] ram_w8_l4096_id7_0_0_rdata,
  input [8-1:0] ram_w8_l4096_id7_0_0_wdata,
  input ram_w8_l4096_id7_0_0_wenable,
  input ram_w8_l4096_id7_0_0_enable,
  input [10-1:0] ram_w8_l4096_id7_0_1_addr,
  output [8-1:0] ram_w8_l4096_id7_0_1_rdata,
  input [8-1:0] ram_w8_l4096_id7_0_1_wdata,
  input ram_w8_l4096_id7_0_1_wenable,
  input ram_w8_l4096_id7_0_1_enable
);

  reg [8-1:0] ram_w8_l4096_id7_0_0_rdata_out;
  assign ram_w8_l4096_id7_0_0_rdata = ram_w8_l4096_id7_0_0_rdata_out;
  reg [8-1:0] ram_w8_l4096_id7_0_1_rdata_out;
  assign ram_w8_l4096_id7_0_1_rdata = ram_w8_l4096_id7_0_1_rdata_out;
  reg [8-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w8_l4096_id7_0_0_enable) begin
      if(ram_w8_l4096_id7_0_0_wenable) begin
        mem[ram_w8_l4096_id7_0_0_addr] <= ram_w8_l4096_id7_0_0_wdata;
        ram_w8_l4096_id7_0_0_rdata_out <= ram_w8_l4096_id7_0_0_wdata;
      end else begin
        ram_w8_l4096_id7_0_0_rdata_out <= mem[ram_w8_l4096_id7_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l4096_id7_0_1_enable) begin
      if(ram_w8_l4096_id7_0_1_wenable) begin
        mem[ram_w8_l4096_id7_0_1_addr] <= ram_w8_l4096_id7_0_1_wdata;
        ram_w8_l4096_id7_0_1_rdata_out <= ram_w8_l4096_id7_0_1_wdata;
      end else begin
        ram_w8_l4096_id7_0_1_rdata_out <= mem[ram_w8_l4096_id7_0_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l4096_id7_1
(
  input CLK,
  input [10-1:0] ram_w8_l4096_id7_1_0_addr,
  output [8-1:0] ram_w8_l4096_id7_1_0_rdata,
  input [8-1:0] ram_w8_l4096_id7_1_0_wdata,
  input ram_w8_l4096_id7_1_0_wenable,
  input ram_w8_l4096_id7_1_0_enable,
  input [10-1:0] ram_w8_l4096_id7_1_1_addr,
  output [8-1:0] ram_w8_l4096_id7_1_1_rdata,
  input [8-1:0] ram_w8_l4096_id7_1_1_wdata,
  input ram_w8_l4096_id7_1_1_wenable,
  input ram_w8_l4096_id7_1_1_enable
);

  reg [8-1:0] ram_w8_l4096_id7_1_0_rdata_out;
  assign ram_w8_l4096_id7_1_0_rdata = ram_w8_l4096_id7_1_0_rdata_out;
  reg [8-1:0] ram_w8_l4096_id7_1_1_rdata_out;
  assign ram_w8_l4096_id7_1_1_rdata = ram_w8_l4096_id7_1_1_rdata_out;
  reg [8-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w8_l4096_id7_1_0_enable) begin
      if(ram_w8_l4096_id7_1_0_wenable) begin
        mem[ram_w8_l4096_id7_1_0_addr] <= ram_w8_l4096_id7_1_0_wdata;
        ram_w8_l4096_id7_1_0_rdata_out <= ram_w8_l4096_id7_1_0_wdata;
      end else begin
        ram_w8_l4096_id7_1_0_rdata_out <= mem[ram_w8_l4096_id7_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l4096_id7_1_1_enable) begin
      if(ram_w8_l4096_id7_1_1_wenable) begin
        mem[ram_w8_l4096_id7_1_1_addr] <= ram_w8_l4096_id7_1_1_wdata;
        ram_w8_l4096_id7_1_1_rdata_out <= ram_w8_l4096_id7_1_1_wdata;
      end else begin
        ram_w8_l4096_id7_1_1_rdata_out <= mem[ram_w8_l4096_id7_1_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l4096_id7_2
(
  input CLK,
  input [10-1:0] ram_w8_l4096_id7_2_0_addr,
  output [8-1:0] ram_w8_l4096_id7_2_0_rdata,
  input [8-1:0] ram_w8_l4096_id7_2_0_wdata,
  input ram_w8_l4096_id7_2_0_wenable,
  input ram_w8_l4096_id7_2_0_enable,
  input [10-1:0] ram_w8_l4096_id7_2_1_addr,
  output [8-1:0] ram_w8_l4096_id7_2_1_rdata,
  input [8-1:0] ram_w8_l4096_id7_2_1_wdata,
  input ram_w8_l4096_id7_2_1_wenable,
  input ram_w8_l4096_id7_2_1_enable
);

  reg [8-1:0] ram_w8_l4096_id7_2_0_rdata_out;
  assign ram_w8_l4096_id7_2_0_rdata = ram_w8_l4096_id7_2_0_rdata_out;
  reg [8-1:0] ram_w8_l4096_id7_2_1_rdata_out;
  assign ram_w8_l4096_id7_2_1_rdata = ram_w8_l4096_id7_2_1_rdata_out;
  reg [8-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w8_l4096_id7_2_0_enable) begin
      if(ram_w8_l4096_id7_2_0_wenable) begin
        mem[ram_w8_l4096_id7_2_0_addr] <= ram_w8_l4096_id7_2_0_wdata;
        ram_w8_l4096_id7_2_0_rdata_out <= ram_w8_l4096_id7_2_0_wdata;
      end else begin
        ram_w8_l4096_id7_2_0_rdata_out <= mem[ram_w8_l4096_id7_2_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l4096_id7_2_1_enable) begin
      if(ram_w8_l4096_id7_2_1_wenable) begin
        mem[ram_w8_l4096_id7_2_1_addr] <= ram_w8_l4096_id7_2_1_wdata;
        ram_w8_l4096_id7_2_1_rdata_out <= ram_w8_l4096_id7_2_1_wdata;
      end else begin
        ram_w8_l4096_id7_2_1_rdata_out <= mem[ram_w8_l4096_id7_2_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l4096_id7_3
(
  input CLK,
  input [10-1:0] ram_w8_l4096_id7_3_0_addr,
  output [8-1:0] ram_w8_l4096_id7_3_0_rdata,
  input [8-1:0] ram_w8_l4096_id7_3_0_wdata,
  input ram_w8_l4096_id7_3_0_wenable,
  input ram_w8_l4096_id7_3_0_enable,
  input [10-1:0] ram_w8_l4096_id7_3_1_addr,
  output [8-1:0] ram_w8_l4096_id7_3_1_rdata,
  input [8-1:0] ram_w8_l4096_id7_3_1_wdata,
  input ram_w8_l4096_id7_3_1_wenable,
  input ram_w8_l4096_id7_3_1_enable
);

  reg [8-1:0] ram_w8_l4096_id7_3_0_rdata_out;
  assign ram_w8_l4096_id7_3_0_rdata = ram_w8_l4096_id7_3_0_rdata_out;
  reg [8-1:0] ram_w8_l4096_id7_3_1_rdata_out;
  assign ram_w8_l4096_id7_3_1_rdata = ram_w8_l4096_id7_3_1_rdata_out;
  reg [8-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w8_l4096_id7_3_0_enable) begin
      if(ram_w8_l4096_id7_3_0_wenable) begin
        mem[ram_w8_l4096_id7_3_0_addr] <= ram_w8_l4096_id7_3_0_wdata;
        ram_w8_l4096_id7_3_0_rdata_out <= ram_w8_l4096_id7_3_0_wdata;
      end else begin
        ram_w8_l4096_id7_3_0_rdata_out <= mem[ram_w8_l4096_id7_3_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l4096_id7_3_1_enable) begin
      if(ram_w8_l4096_id7_3_1_wenable) begin
        mem[ram_w8_l4096_id7_3_1_addr] <= ram_w8_l4096_id7_3_1_wdata;
        ram_w8_l4096_id7_3_1_rdata_out <= ram_w8_l4096_id7_3_1_wdata;
      end else begin
        ram_w8_l4096_id7_3_1_rdata_out <= mem[ram_w8_l4096_id7_3_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l4096_id8_0
(
  input CLK,
  input [10-1:0] ram_w8_l4096_id8_0_0_addr,
  output [8-1:0] ram_w8_l4096_id8_0_0_rdata,
  input [8-1:0] ram_w8_l4096_id8_0_0_wdata,
  input ram_w8_l4096_id8_0_0_wenable,
  input ram_w8_l4096_id8_0_0_enable,
  input [10-1:0] ram_w8_l4096_id8_0_1_addr,
  output [8-1:0] ram_w8_l4096_id8_0_1_rdata,
  input [8-1:0] ram_w8_l4096_id8_0_1_wdata,
  input ram_w8_l4096_id8_0_1_wenable,
  input ram_w8_l4096_id8_0_1_enable
);

  reg [8-1:0] ram_w8_l4096_id8_0_0_rdata_out;
  assign ram_w8_l4096_id8_0_0_rdata = ram_w8_l4096_id8_0_0_rdata_out;
  reg [8-1:0] ram_w8_l4096_id8_0_1_rdata_out;
  assign ram_w8_l4096_id8_0_1_rdata = ram_w8_l4096_id8_0_1_rdata_out;
  reg [8-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w8_l4096_id8_0_0_enable) begin
      if(ram_w8_l4096_id8_0_0_wenable) begin
        mem[ram_w8_l4096_id8_0_0_addr] <= ram_w8_l4096_id8_0_0_wdata;
        ram_w8_l4096_id8_0_0_rdata_out <= ram_w8_l4096_id8_0_0_wdata;
      end else begin
        ram_w8_l4096_id8_0_0_rdata_out <= mem[ram_w8_l4096_id8_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l4096_id8_0_1_enable) begin
      if(ram_w8_l4096_id8_0_1_wenable) begin
        mem[ram_w8_l4096_id8_0_1_addr] <= ram_w8_l4096_id8_0_1_wdata;
        ram_w8_l4096_id8_0_1_rdata_out <= ram_w8_l4096_id8_0_1_wdata;
      end else begin
        ram_w8_l4096_id8_0_1_rdata_out <= mem[ram_w8_l4096_id8_0_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l4096_id8_1
(
  input CLK,
  input [10-1:0] ram_w8_l4096_id8_1_0_addr,
  output [8-1:0] ram_w8_l4096_id8_1_0_rdata,
  input [8-1:0] ram_w8_l4096_id8_1_0_wdata,
  input ram_w8_l4096_id8_1_0_wenable,
  input ram_w8_l4096_id8_1_0_enable,
  input [10-1:0] ram_w8_l4096_id8_1_1_addr,
  output [8-1:0] ram_w8_l4096_id8_1_1_rdata,
  input [8-1:0] ram_w8_l4096_id8_1_1_wdata,
  input ram_w8_l4096_id8_1_1_wenable,
  input ram_w8_l4096_id8_1_1_enable
);

  reg [8-1:0] ram_w8_l4096_id8_1_0_rdata_out;
  assign ram_w8_l4096_id8_1_0_rdata = ram_w8_l4096_id8_1_0_rdata_out;
  reg [8-1:0] ram_w8_l4096_id8_1_1_rdata_out;
  assign ram_w8_l4096_id8_1_1_rdata = ram_w8_l4096_id8_1_1_rdata_out;
  reg [8-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w8_l4096_id8_1_0_enable) begin
      if(ram_w8_l4096_id8_1_0_wenable) begin
        mem[ram_w8_l4096_id8_1_0_addr] <= ram_w8_l4096_id8_1_0_wdata;
        ram_w8_l4096_id8_1_0_rdata_out <= ram_w8_l4096_id8_1_0_wdata;
      end else begin
        ram_w8_l4096_id8_1_0_rdata_out <= mem[ram_w8_l4096_id8_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l4096_id8_1_1_enable) begin
      if(ram_w8_l4096_id8_1_1_wenable) begin
        mem[ram_w8_l4096_id8_1_1_addr] <= ram_w8_l4096_id8_1_1_wdata;
        ram_w8_l4096_id8_1_1_rdata_out <= ram_w8_l4096_id8_1_1_wdata;
      end else begin
        ram_w8_l4096_id8_1_1_rdata_out <= mem[ram_w8_l4096_id8_1_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l4096_id8_2
(
  input CLK,
  input [10-1:0] ram_w8_l4096_id8_2_0_addr,
  output [8-1:0] ram_w8_l4096_id8_2_0_rdata,
  input [8-1:0] ram_w8_l4096_id8_2_0_wdata,
  input ram_w8_l4096_id8_2_0_wenable,
  input ram_w8_l4096_id8_2_0_enable,
  input [10-1:0] ram_w8_l4096_id8_2_1_addr,
  output [8-1:0] ram_w8_l4096_id8_2_1_rdata,
  input [8-1:0] ram_w8_l4096_id8_2_1_wdata,
  input ram_w8_l4096_id8_2_1_wenable,
  input ram_w8_l4096_id8_2_1_enable
);

  reg [8-1:0] ram_w8_l4096_id8_2_0_rdata_out;
  assign ram_w8_l4096_id8_2_0_rdata = ram_w8_l4096_id8_2_0_rdata_out;
  reg [8-1:0] ram_w8_l4096_id8_2_1_rdata_out;
  assign ram_w8_l4096_id8_2_1_rdata = ram_w8_l4096_id8_2_1_rdata_out;
  reg [8-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w8_l4096_id8_2_0_enable) begin
      if(ram_w8_l4096_id8_2_0_wenable) begin
        mem[ram_w8_l4096_id8_2_0_addr] <= ram_w8_l4096_id8_2_0_wdata;
        ram_w8_l4096_id8_2_0_rdata_out <= ram_w8_l4096_id8_2_0_wdata;
      end else begin
        ram_w8_l4096_id8_2_0_rdata_out <= mem[ram_w8_l4096_id8_2_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l4096_id8_2_1_enable) begin
      if(ram_w8_l4096_id8_2_1_wenable) begin
        mem[ram_w8_l4096_id8_2_1_addr] <= ram_w8_l4096_id8_2_1_wdata;
        ram_w8_l4096_id8_2_1_rdata_out <= ram_w8_l4096_id8_2_1_wdata;
      end else begin
        ram_w8_l4096_id8_2_1_rdata_out <= mem[ram_w8_l4096_id8_2_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l4096_id8_3
(
  input CLK,
  input [10-1:0] ram_w8_l4096_id8_3_0_addr,
  output [8-1:0] ram_w8_l4096_id8_3_0_rdata,
  input [8-1:0] ram_w8_l4096_id8_3_0_wdata,
  input ram_w8_l4096_id8_3_0_wenable,
  input ram_w8_l4096_id8_3_0_enable,
  input [10-1:0] ram_w8_l4096_id8_3_1_addr,
  output [8-1:0] ram_w8_l4096_id8_3_1_rdata,
  input [8-1:0] ram_w8_l4096_id8_3_1_wdata,
  input ram_w8_l4096_id8_3_1_wenable,
  input ram_w8_l4096_id8_3_1_enable
);

  reg [8-1:0] ram_w8_l4096_id8_3_0_rdata_out;
  assign ram_w8_l4096_id8_3_0_rdata = ram_w8_l4096_id8_3_0_rdata_out;
  reg [8-1:0] ram_w8_l4096_id8_3_1_rdata_out;
  assign ram_w8_l4096_id8_3_1_rdata = ram_w8_l4096_id8_3_1_rdata_out;
  reg [8-1:0] mem [0:1024-1];

  always @(posedge CLK) begin
    if(ram_w8_l4096_id8_3_0_enable) begin
      if(ram_w8_l4096_id8_3_0_wenable) begin
        mem[ram_w8_l4096_id8_3_0_addr] <= ram_w8_l4096_id8_3_0_wdata;
        ram_w8_l4096_id8_3_0_rdata_out <= ram_w8_l4096_id8_3_0_wdata;
      end else begin
        ram_w8_l4096_id8_3_0_rdata_out <= mem[ram_w8_l4096_id8_3_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l4096_id8_3_1_enable) begin
      if(ram_w8_l4096_id8_3_1_wenable) begin
        mem[ram_w8_l4096_id8_3_1_addr] <= ram_w8_l4096_id8_3_1_wdata;
        ram_w8_l4096_id8_3_1_rdata_out <= ram_w8_l4096_id8_3_1_wdata;
      end else begin
        ram_w8_l4096_id8_3_1_rdata_out <= mem[ram_w8_l4096_id8_3_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l2048_id0_0
(
  input CLK,
  input [9-1:0] ram_w8_l2048_id0_0_0_addr,
  output [8-1:0] ram_w8_l2048_id0_0_0_rdata,
  input [8-1:0] ram_w8_l2048_id0_0_0_wdata,
  input ram_w8_l2048_id0_0_0_wenable,
  input ram_w8_l2048_id0_0_0_enable,
  input [9-1:0] ram_w8_l2048_id0_0_1_addr,
  output [8-1:0] ram_w8_l2048_id0_0_1_rdata,
  input [8-1:0] ram_w8_l2048_id0_0_1_wdata,
  input ram_w8_l2048_id0_0_1_wenable,
  input ram_w8_l2048_id0_0_1_enable
);

  reg [8-1:0] ram_w8_l2048_id0_0_0_rdata_out;
  assign ram_w8_l2048_id0_0_0_rdata = ram_w8_l2048_id0_0_0_rdata_out;
  reg [8-1:0] ram_w8_l2048_id0_0_1_rdata_out;
  assign ram_w8_l2048_id0_0_1_rdata = ram_w8_l2048_id0_0_1_rdata_out;
  reg [8-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id0_0_0_enable) begin
      if(ram_w8_l2048_id0_0_0_wenable) begin
        mem[ram_w8_l2048_id0_0_0_addr] <= ram_w8_l2048_id0_0_0_wdata;
        ram_w8_l2048_id0_0_0_rdata_out <= ram_w8_l2048_id0_0_0_wdata;
      end else begin
        ram_w8_l2048_id0_0_0_rdata_out <= mem[ram_w8_l2048_id0_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l2048_id0_0_1_enable) begin
      if(ram_w8_l2048_id0_0_1_wenable) begin
        mem[ram_w8_l2048_id0_0_1_addr] <= ram_w8_l2048_id0_0_1_wdata;
        ram_w8_l2048_id0_0_1_rdata_out <= ram_w8_l2048_id0_0_1_wdata;
      end else begin
        ram_w8_l2048_id0_0_1_rdata_out <= mem[ram_w8_l2048_id0_0_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l2048_id0_1
(
  input CLK,
  input [9-1:0] ram_w8_l2048_id0_1_0_addr,
  output [8-1:0] ram_w8_l2048_id0_1_0_rdata,
  input [8-1:0] ram_w8_l2048_id0_1_0_wdata,
  input ram_w8_l2048_id0_1_0_wenable,
  input ram_w8_l2048_id0_1_0_enable,
  input [9-1:0] ram_w8_l2048_id0_1_1_addr,
  output [8-1:0] ram_w8_l2048_id0_1_1_rdata,
  input [8-1:0] ram_w8_l2048_id0_1_1_wdata,
  input ram_w8_l2048_id0_1_1_wenable,
  input ram_w8_l2048_id0_1_1_enable
);

  reg [8-1:0] ram_w8_l2048_id0_1_0_rdata_out;
  assign ram_w8_l2048_id0_1_0_rdata = ram_w8_l2048_id0_1_0_rdata_out;
  reg [8-1:0] ram_w8_l2048_id0_1_1_rdata_out;
  assign ram_w8_l2048_id0_1_1_rdata = ram_w8_l2048_id0_1_1_rdata_out;
  reg [8-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id0_1_0_enable) begin
      if(ram_w8_l2048_id0_1_0_wenable) begin
        mem[ram_w8_l2048_id0_1_0_addr] <= ram_w8_l2048_id0_1_0_wdata;
        ram_w8_l2048_id0_1_0_rdata_out <= ram_w8_l2048_id0_1_0_wdata;
      end else begin
        ram_w8_l2048_id0_1_0_rdata_out <= mem[ram_w8_l2048_id0_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l2048_id0_1_1_enable) begin
      if(ram_w8_l2048_id0_1_1_wenable) begin
        mem[ram_w8_l2048_id0_1_1_addr] <= ram_w8_l2048_id0_1_1_wdata;
        ram_w8_l2048_id0_1_1_rdata_out <= ram_w8_l2048_id0_1_1_wdata;
      end else begin
        ram_w8_l2048_id0_1_1_rdata_out <= mem[ram_w8_l2048_id0_1_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l2048_id0_2
(
  input CLK,
  input [9-1:0] ram_w8_l2048_id0_2_0_addr,
  output [8-1:0] ram_w8_l2048_id0_2_0_rdata,
  input [8-1:0] ram_w8_l2048_id0_2_0_wdata,
  input ram_w8_l2048_id0_2_0_wenable,
  input ram_w8_l2048_id0_2_0_enable,
  input [9-1:0] ram_w8_l2048_id0_2_1_addr,
  output [8-1:0] ram_w8_l2048_id0_2_1_rdata,
  input [8-1:0] ram_w8_l2048_id0_2_1_wdata,
  input ram_w8_l2048_id0_2_1_wenable,
  input ram_w8_l2048_id0_2_1_enable
);

  reg [8-1:0] ram_w8_l2048_id0_2_0_rdata_out;
  assign ram_w8_l2048_id0_2_0_rdata = ram_w8_l2048_id0_2_0_rdata_out;
  reg [8-1:0] ram_w8_l2048_id0_2_1_rdata_out;
  assign ram_w8_l2048_id0_2_1_rdata = ram_w8_l2048_id0_2_1_rdata_out;
  reg [8-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id0_2_0_enable) begin
      if(ram_w8_l2048_id0_2_0_wenable) begin
        mem[ram_w8_l2048_id0_2_0_addr] <= ram_w8_l2048_id0_2_0_wdata;
        ram_w8_l2048_id0_2_0_rdata_out <= ram_w8_l2048_id0_2_0_wdata;
      end else begin
        ram_w8_l2048_id0_2_0_rdata_out <= mem[ram_w8_l2048_id0_2_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l2048_id0_2_1_enable) begin
      if(ram_w8_l2048_id0_2_1_wenable) begin
        mem[ram_w8_l2048_id0_2_1_addr] <= ram_w8_l2048_id0_2_1_wdata;
        ram_w8_l2048_id0_2_1_rdata_out <= ram_w8_l2048_id0_2_1_wdata;
      end else begin
        ram_w8_l2048_id0_2_1_rdata_out <= mem[ram_w8_l2048_id0_2_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l2048_id0_3
(
  input CLK,
  input [9-1:0] ram_w8_l2048_id0_3_0_addr,
  output [8-1:0] ram_w8_l2048_id0_3_0_rdata,
  input [8-1:0] ram_w8_l2048_id0_3_0_wdata,
  input ram_w8_l2048_id0_3_0_wenable,
  input ram_w8_l2048_id0_3_0_enable,
  input [9-1:0] ram_w8_l2048_id0_3_1_addr,
  output [8-1:0] ram_w8_l2048_id0_3_1_rdata,
  input [8-1:0] ram_w8_l2048_id0_3_1_wdata,
  input ram_w8_l2048_id0_3_1_wenable,
  input ram_w8_l2048_id0_3_1_enable
);

  reg [8-1:0] ram_w8_l2048_id0_3_0_rdata_out;
  assign ram_w8_l2048_id0_3_0_rdata = ram_w8_l2048_id0_3_0_rdata_out;
  reg [8-1:0] ram_w8_l2048_id0_3_1_rdata_out;
  assign ram_w8_l2048_id0_3_1_rdata = ram_w8_l2048_id0_3_1_rdata_out;
  reg [8-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id0_3_0_enable) begin
      if(ram_w8_l2048_id0_3_0_wenable) begin
        mem[ram_w8_l2048_id0_3_0_addr] <= ram_w8_l2048_id0_3_0_wdata;
        ram_w8_l2048_id0_3_0_rdata_out <= ram_w8_l2048_id0_3_0_wdata;
      end else begin
        ram_w8_l2048_id0_3_0_rdata_out <= mem[ram_w8_l2048_id0_3_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l2048_id0_3_1_enable) begin
      if(ram_w8_l2048_id0_3_1_wenable) begin
        mem[ram_w8_l2048_id0_3_1_addr] <= ram_w8_l2048_id0_3_1_wdata;
        ram_w8_l2048_id0_3_1_rdata_out <= ram_w8_l2048_id0_3_1_wdata;
      end else begin
        ram_w8_l2048_id0_3_1_rdata_out <= mem[ram_w8_l2048_id0_3_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l2048_id1_0
(
  input CLK,
  input [9-1:0] ram_w8_l2048_id1_0_0_addr,
  output [8-1:0] ram_w8_l2048_id1_0_0_rdata,
  input [8-1:0] ram_w8_l2048_id1_0_0_wdata,
  input ram_w8_l2048_id1_0_0_wenable,
  input ram_w8_l2048_id1_0_0_enable,
  input [9-1:0] ram_w8_l2048_id1_0_1_addr,
  output [8-1:0] ram_w8_l2048_id1_0_1_rdata,
  input [8-1:0] ram_w8_l2048_id1_0_1_wdata,
  input ram_w8_l2048_id1_0_1_wenable,
  input ram_w8_l2048_id1_0_1_enable
);

  reg [8-1:0] ram_w8_l2048_id1_0_0_rdata_out;
  assign ram_w8_l2048_id1_0_0_rdata = ram_w8_l2048_id1_0_0_rdata_out;
  reg [8-1:0] ram_w8_l2048_id1_0_1_rdata_out;
  assign ram_w8_l2048_id1_0_1_rdata = ram_w8_l2048_id1_0_1_rdata_out;
  reg [8-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id1_0_0_enable) begin
      if(ram_w8_l2048_id1_0_0_wenable) begin
        mem[ram_w8_l2048_id1_0_0_addr] <= ram_w8_l2048_id1_0_0_wdata;
        ram_w8_l2048_id1_0_0_rdata_out <= ram_w8_l2048_id1_0_0_wdata;
      end else begin
        ram_w8_l2048_id1_0_0_rdata_out <= mem[ram_w8_l2048_id1_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l2048_id1_0_1_enable) begin
      if(ram_w8_l2048_id1_0_1_wenable) begin
        mem[ram_w8_l2048_id1_0_1_addr] <= ram_w8_l2048_id1_0_1_wdata;
        ram_w8_l2048_id1_0_1_rdata_out <= ram_w8_l2048_id1_0_1_wdata;
      end else begin
        ram_w8_l2048_id1_0_1_rdata_out <= mem[ram_w8_l2048_id1_0_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l2048_id1_1
(
  input CLK,
  input [9-1:0] ram_w8_l2048_id1_1_0_addr,
  output [8-1:0] ram_w8_l2048_id1_1_0_rdata,
  input [8-1:0] ram_w8_l2048_id1_1_0_wdata,
  input ram_w8_l2048_id1_1_0_wenable,
  input ram_w8_l2048_id1_1_0_enable,
  input [9-1:0] ram_w8_l2048_id1_1_1_addr,
  output [8-1:0] ram_w8_l2048_id1_1_1_rdata,
  input [8-1:0] ram_w8_l2048_id1_1_1_wdata,
  input ram_w8_l2048_id1_1_1_wenable,
  input ram_w8_l2048_id1_1_1_enable
);

  reg [8-1:0] ram_w8_l2048_id1_1_0_rdata_out;
  assign ram_w8_l2048_id1_1_0_rdata = ram_w8_l2048_id1_1_0_rdata_out;
  reg [8-1:0] ram_w8_l2048_id1_1_1_rdata_out;
  assign ram_w8_l2048_id1_1_1_rdata = ram_w8_l2048_id1_1_1_rdata_out;
  reg [8-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id1_1_0_enable) begin
      if(ram_w8_l2048_id1_1_0_wenable) begin
        mem[ram_w8_l2048_id1_1_0_addr] <= ram_w8_l2048_id1_1_0_wdata;
        ram_w8_l2048_id1_1_0_rdata_out <= ram_w8_l2048_id1_1_0_wdata;
      end else begin
        ram_w8_l2048_id1_1_0_rdata_out <= mem[ram_w8_l2048_id1_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l2048_id1_1_1_enable) begin
      if(ram_w8_l2048_id1_1_1_wenable) begin
        mem[ram_w8_l2048_id1_1_1_addr] <= ram_w8_l2048_id1_1_1_wdata;
        ram_w8_l2048_id1_1_1_rdata_out <= ram_w8_l2048_id1_1_1_wdata;
      end else begin
        ram_w8_l2048_id1_1_1_rdata_out <= mem[ram_w8_l2048_id1_1_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l2048_id1_2
(
  input CLK,
  input [9-1:0] ram_w8_l2048_id1_2_0_addr,
  output [8-1:0] ram_w8_l2048_id1_2_0_rdata,
  input [8-1:0] ram_w8_l2048_id1_2_0_wdata,
  input ram_w8_l2048_id1_2_0_wenable,
  input ram_w8_l2048_id1_2_0_enable,
  input [9-1:0] ram_w8_l2048_id1_2_1_addr,
  output [8-1:0] ram_w8_l2048_id1_2_1_rdata,
  input [8-1:0] ram_w8_l2048_id1_2_1_wdata,
  input ram_w8_l2048_id1_2_1_wenable,
  input ram_w8_l2048_id1_2_1_enable
);

  reg [8-1:0] ram_w8_l2048_id1_2_0_rdata_out;
  assign ram_w8_l2048_id1_2_0_rdata = ram_w8_l2048_id1_2_0_rdata_out;
  reg [8-1:0] ram_w8_l2048_id1_2_1_rdata_out;
  assign ram_w8_l2048_id1_2_1_rdata = ram_w8_l2048_id1_2_1_rdata_out;
  reg [8-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id1_2_0_enable) begin
      if(ram_w8_l2048_id1_2_0_wenable) begin
        mem[ram_w8_l2048_id1_2_0_addr] <= ram_w8_l2048_id1_2_0_wdata;
        ram_w8_l2048_id1_2_0_rdata_out <= ram_w8_l2048_id1_2_0_wdata;
      end else begin
        ram_w8_l2048_id1_2_0_rdata_out <= mem[ram_w8_l2048_id1_2_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l2048_id1_2_1_enable) begin
      if(ram_w8_l2048_id1_2_1_wenable) begin
        mem[ram_w8_l2048_id1_2_1_addr] <= ram_w8_l2048_id1_2_1_wdata;
        ram_w8_l2048_id1_2_1_rdata_out <= ram_w8_l2048_id1_2_1_wdata;
      end else begin
        ram_w8_l2048_id1_2_1_rdata_out <= mem[ram_w8_l2048_id1_2_1_addr];
      end
    end 
  end


endmodule



module ram_w8_l2048_id1_3
(
  input CLK,
  input [9-1:0] ram_w8_l2048_id1_3_0_addr,
  output [8-1:0] ram_w8_l2048_id1_3_0_rdata,
  input [8-1:0] ram_w8_l2048_id1_3_0_wdata,
  input ram_w8_l2048_id1_3_0_wenable,
  input ram_w8_l2048_id1_3_0_enable,
  input [9-1:0] ram_w8_l2048_id1_3_1_addr,
  output [8-1:0] ram_w8_l2048_id1_3_1_rdata,
  input [8-1:0] ram_w8_l2048_id1_3_1_wdata,
  input ram_w8_l2048_id1_3_1_wenable,
  input ram_w8_l2048_id1_3_1_enable
);

  reg [8-1:0] ram_w8_l2048_id1_3_0_rdata_out;
  assign ram_w8_l2048_id1_3_0_rdata = ram_w8_l2048_id1_3_0_rdata_out;
  reg [8-1:0] ram_w8_l2048_id1_3_1_rdata_out;
  assign ram_w8_l2048_id1_3_1_rdata = ram_w8_l2048_id1_3_1_rdata_out;
  reg [8-1:0] mem [0:512-1];

  always @(posedge CLK) begin
    if(ram_w8_l2048_id1_3_0_enable) begin
      if(ram_w8_l2048_id1_3_0_wenable) begin
        mem[ram_w8_l2048_id1_3_0_addr] <= ram_w8_l2048_id1_3_0_wdata;
        ram_w8_l2048_id1_3_0_rdata_out <= ram_w8_l2048_id1_3_0_wdata;
      end else begin
        ram_w8_l2048_id1_3_0_rdata_out <= mem[ram_w8_l2048_id1_3_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w8_l2048_id1_3_1_enable) begin
      if(ram_w8_l2048_id1_3_1_wenable) begin
        mem[ram_w8_l2048_id1_3_1_addr] <= ram_w8_l2048_id1_3_1_wdata;
        ram_w8_l2048_id1_3_1_rdata_out <= ram_w8_l2048_id1_3_1_wdata;
      end else begin
        ram_w8_l2048_id1_3_1_rdata_out <= mem[ram_w8_l2048_id1_3_1_addr];
      end
    end 
  end


endmodule



module madd_0
(
  input CLK,
  input update,
  input [8-1:0] a,
  input [8-1:0] b,
  input [8-1:0] c,
  output [16-1:0] d
);


  madd_core_0
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_0
(
  input CLK,
  input update,
  input [8-1:0] a,
  input [8-1:0] b,
  input [8-1:0] c,
  output [16-1:0] d
);

  reg signed [8-1:0] _a;
  reg signed [8-1:0] _b;
  reg signed [8-1:0] _c;
  wire signed [16-1:0] _mul;
  wire signed [16-1:0] _madd;
  reg signed [16-1:0] _pipe_madd0;
  reg signed [16-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_1
(
  input CLK,
  input update,
  input [8-1:0] a,
  input [8-1:0] b,
  input [8-1:0] c,
  output [16-1:0] d
);


  madd_core_1
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_1
(
  input CLK,
  input update,
  input [8-1:0] a,
  input [8-1:0] b,
  input [8-1:0] c,
  output [16-1:0] d
);

  reg signed [8-1:0] _a;
  reg signed [8-1:0] _b;
  reg signed [8-1:0] _c;
  wire signed [16-1:0] _mul;
  wire signed [16-1:0] _madd;
  reg signed [16-1:0] _pipe_madd0;
  reg signed [16-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_2
(
  input CLK,
  input update,
  input [8-1:0] a,
  input [8-1:0] b,
  input [8-1:0] c,
  output [16-1:0] d
);


  madd_core_2
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_2
(
  input CLK,
  input update,
  input [8-1:0] a,
  input [8-1:0] b,
  input [8-1:0] c,
  output [16-1:0] d
);

  reg signed [8-1:0] _a;
  reg signed [8-1:0] _b;
  reg signed [8-1:0] _c;
  wire signed [16-1:0] _mul;
  wire signed [16-1:0] _madd;
  reg signed [16-1:0] _pipe_madd0;
  reg signed [16-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_3
(
  input CLK,
  input update,
  input [8-1:0] a,
  input [8-1:0] b,
  input [8-1:0] c,
  output [16-1:0] d
);


  madd_core_3
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_3
(
  input CLK,
  input update,
  input [8-1:0] a,
  input [8-1:0] b,
  input [8-1:0] c,
  output [16-1:0] d
);

  reg signed [8-1:0] _a;
  reg signed [8-1:0] _b;
  reg signed [8-1:0] _c;
  wire signed [16-1:0] _mul;
  wire signed [16-1:0] _madd;
  reg signed [16-1:0] _pipe_madd0;
  reg signed [16-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_4
(
  input CLK,
  input update,
  input [8-1:0] a,
  input [8-1:0] b,
  input [8-1:0] c,
  output [16-1:0] d
);


  madd_core_4
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_4
(
  input CLK,
  input update,
  input [8-1:0] a,
  input [8-1:0] b,
  input [8-1:0] c,
  output [16-1:0] d
);

  reg signed [8-1:0] _a;
  reg signed [8-1:0] _b;
  reg signed [8-1:0] _c;
  wire signed [16-1:0] _mul;
  wire signed [16-1:0] _madd;
  reg signed [16-1:0] _pipe_madd0;
  reg signed [16-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_5
(
  input CLK,
  input update,
  input [8-1:0] a,
  input [8-1:0] b,
  input [8-1:0] c,
  output [16-1:0] d
);


  madd_core_5
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_5
(
  input CLK,
  input update,
  input [8-1:0] a,
  input [8-1:0] b,
  input [8-1:0] c,
  output [16-1:0] d
);

  reg signed [8-1:0] _a;
  reg signed [8-1:0] _b;
  reg signed [8-1:0] _c;
  wire signed [16-1:0] _mul;
  wire signed [16-1:0] _madd;
  reg signed [16-1:0] _pipe_madd0;
  reg signed [16-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_6
(
  input CLK,
  input update,
  input [8-1:0] a,
  input [8-1:0] b,
  input [8-1:0] c,
  output [16-1:0] d
);


  madd_core_6
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_6
(
  input CLK,
  input update,
  input [8-1:0] a,
  input [8-1:0] b,
  input [8-1:0] c,
  output [16-1:0] d
);

  reg signed [8-1:0] _a;
  reg signed [8-1:0] _b;
  reg signed [8-1:0] _c;
  wire signed [16-1:0] _mul;
  wire signed [16-1:0] _madd;
  reg signed [16-1:0] _pipe_madd0;
  reg signed [16-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_7
(
  input CLK,
  input update,
  input [8-1:0] a,
  input [8-1:0] b,
  input [8-1:0] c,
  output [16-1:0] d
);


  madd_core_7
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_7
(
  input CLK,
  input update,
  input [8-1:0] a,
  input [8-1:0] b,
  input [8-1:0] c,
  output [16-1:0] d
);

  reg signed [8-1:0] _a;
  reg signed [8-1:0] _b;
  reg signed [8-1:0] _c;
  wire signed [16-1:0] _mul;
  wire signed [16-1:0] _madd;
  reg signed [16-1:0] _pipe_madd0;
  reg signed [16-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_8
(
  input CLK,
  input update,
  input [8-1:0] a,
  input [8-1:0] b,
  input [8-1:0] c,
  output [16-1:0] d
);


  madd_core_8
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_8
(
  input CLK,
  input update,
  input [8-1:0] a,
  input [8-1:0] b,
  input [8-1:0] c,
  output [16-1:0] d
);

  reg signed [8-1:0] _a;
  reg signed [8-1:0] _b;
  reg signed [8-1:0] _c;
  wire signed [16-1:0] _mul;
  wire signed [16-1:0] _madd;
  reg signed [16-1:0] _pipe_madd0;
  reg signed [16-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module multiplier_0
(
  input CLK,
  input update,
  input [32-1:0] a,
  input [8-1:0] b,
  output [40-1:0] c
);


  multiplier_core_0
  mult
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c)
  );


endmodule



module multiplier_core_0
(
  input CLK,
  input update,
  input [32-1:0] a,
  input [8-1:0] b,
  output [40-1:0] c
);

  reg signed [32-1:0] _a;
  reg signed [8-1:0] _b;
  wire signed [40-1:0] _mul;
  reg signed [40-1:0] _pipe_mul0;
  reg signed [40-1:0] _pipe_mul1;
  assign _mul = _a * _b;
  assign c = _pipe_mul1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _pipe_mul0 <= _mul;
      _pipe_mul1 <= _pipe_mul0;
    end 
  end


endmodule

